../sandbox/bios1_rom-behavior.vhdl