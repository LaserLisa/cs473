../sandbox/bios_rom-entity.vhdl