../sandbox/bios1_rom-entity.vhdl