--------------------------------------------------------------------------------
-- $RCSfile: $
--
-- DESC    : OpenRisk 1420 
--
-- AUTHOR  : Dr. Theo Kluter
--
-- CVS     : $Revision: $
--           $Date: $
--           $Author: $
--           $Source: $
--
--------------------------------------------------------------------------------
--
--  HISTORY :
--
--  $Log: 
--------------------------------------------------------------------------------

ARCHITECTURE platform_independent OF bios_rom IS

BEGIN

   TheRom : PROCESS( address )
   BEGIN
      CASE (address) IS
         WHEN "00000000000" => data <= X"2014ADDE";
         WHEN "00000000001" => data <= X"00000015";
         WHEN "00000000010" => data <= X"11000000";
         WHEN "00000000011" => data <= X"00000015";
         WHEN "00000000100" => data <= X"0F000000";
         WHEN "00000000101" => data <= X"00000015";
         WHEN "00000000110" => data <= X"0D000000";
         WHEN "00000000111" => data <= X"00000015";
         WHEN "00000001000" => data <= X"0B000000";
         WHEN "00000001001" => data <= X"00000015";
         WHEN "00000001010" => data <= X"09000000";
         WHEN "00000001011" => data <= X"00000015";
         WHEN "00000001100" => data <= X"00C02018";
         WHEN "00000001101" => data <= X"FC1F21A8";
         WHEN "00000001110" => data <= X"050060E0";
         WHEN "00000001111" => data <= X"FA020004";
         WHEN "00000010000" => data <= X"050080E0";
         WHEN "00000010010" => data <= X"00000015";
         WHEN "00000010011" => data <= X"84FF219C";
         WHEN "00000010100" => data <= X"001001D4";
         WHEN "00000010101" => data <= X"041801D4";
         WHEN "00000010110" => data <= X"082001D4";
         WHEN "00000010111" => data <= X"0C2801D4";
         WHEN "00000011000" => data <= X"103001D4";
         WHEN "00000011001" => data <= X"143801D4";
         WHEN "00000011010" => data <= X"184001D4";
         WHEN "00000011011" => data <= X"1C4801D4";
         WHEN "00000011100" => data <= X"205001D4";
         WHEN "00000011101" => data <= X"245801D4";
         WHEN "00000011110" => data <= X"286001D4";
         WHEN "00000011111" => data <= X"2C6801D4";
         WHEN "00000100000" => data <= X"307001D4";
         WHEN "00000100001" => data <= X"347801D4";
         WHEN "00000100010" => data <= X"388001D4";
         WHEN "00000100011" => data <= X"3C8801D4";
         WHEN "00000100100" => data <= X"409001D4";
         WHEN "00000100101" => data <= X"449801D4";
         WHEN "00000100110" => data <= X"48A001D4";
         WHEN "00000100111" => data <= X"4CA801D4";
         WHEN "00000101000" => data <= X"50B001D4";
         WHEN "00000101001" => data <= X"54B801D4";
         WHEN "00000101010" => data <= X"58C001D4";
         WHEN "00000101011" => data <= X"5CC801D4";
         WHEN "00000101100" => data <= X"60D001D4";
         WHEN "00000101101" => data <= X"64D801D4";
         WHEN "00000101110" => data <= X"68E001D4";
         WHEN "00000101111" => data <= X"6CE801D4";
         WHEN "00000110000" => data <= X"70F001D4";
         WHEN "00000110001" => data <= X"74F801D4";
         WHEN "00000110010" => data <= X"1200E0B7";
         WHEN "00000110011" => data <= X"0200FFBB";
         WHEN "00000110100" => data <= X"00F0C01B";
         WHEN "00000110101" => data <= X"6C01DEAB";
         WHEN "00000110110" => data <= X"00F8DEE3";
         WHEN "00000110111" => data <= X"0000FE87";
         WHEN "00000111000" => data <= X"00F80048";
         WHEN "00000111001" => data <= X"00000015";
         WHEN "00000111010" => data <= X"00004184";
         WHEN "00000111011" => data <= X"04006184";
         WHEN "00000111100" => data <= X"08008184";
         WHEN "00000111101" => data <= X"0C00A184";
         WHEN "00000111110" => data <= X"1000C184";
         WHEN "00000111111" => data <= X"1400E184";
         WHEN "00001000000" => data <= X"18000185";
         WHEN "00001000001" => data <= X"1C002185";
         WHEN "00001000010" => data <= X"20004185";
         WHEN "00001000011" => data <= X"24006185";
         WHEN "00001000100" => data <= X"28008185";
         WHEN "00001000101" => data <= X"2C00A185";
         WHEN "00001000110" => data <= X"3000C185";
         WHEN "00001000111" => data <= X"3400E185";
         WHEN "00001001000" => data <= X"38000186";
         WHEN "00001001001" => data <= X"3C002186";
         WHEN "00001001010" => data <= X"40004186";
         WHEN "00001001011" => data <= X"44006186";
         WHEN "00001001100" => data <= X"48008186";
         WHEN "00001001101" => data <= X"4C00A186";
         WHEN "00001001110" => data <= X"5000C186";
         WHEN "00001001111" => data <= X"5400E186";
         WHEN "00001010000" => data <= X"58000187";
         WHEN "00001010001" => data <= X"5C002187";
         WHEN "00001010010" => data <= X"60004187";
         WHEN "00001010011" => data <= X"64006187";
         WHEN "00001010100" => data <= X"68008187";
         WHEN "00001010101" => data <= X"6C00A187";
         WHEN "00001010110" => data <= X"7000C187";
         WHEN "00001010111" => data <= X"7400E187";
         WHEN "00001011000" => data <= X"7C00219C";
         WHEN "00001011001" => data <= X"00000024";
         WHEN "00001011010" => data <= X"00000015";
         WHEN "00001011011" => data <= X"300000F0";
         WHEN "00001011100" => data <= X"840100F0";
         WHEN "00001011101" => data <= X"A00100F0";
         WHEN "00001011110" => data <= X"BC0100F0";
         WHEN "00001011111" => data <= X"D80100F0";
         WHEN "00001100000" => data <= X"F40100F0";
         WHEN "00001100001" => data <= X"00F0A018";
         WHEN "00001100010" => data <= X"00F08018";
         WHEN "00001100011" => data <= X"00F06018";
         WHEN "00001100100" => data <= X"D417A59C";
         WHEN "00001100101" => data <= X"5408849C";
         WHEN "00001100110" => data <= X"2C010000";
         WHEN "00001100111" => data <= X"AC09639C";
         WHEN "00001101000" => data <= X"00F0A018";
         WHEN "00001101001" => data <= X"00F08018";
         WHEN "00001101010" => data <= X"00F06018";
         WHEN "00001101011" => data <= X"DF17A59C";
         WHEN "00001101100" => data <= X"5408849C";
         WHEN "00001101101" => data <= X"25010000";
         WHEN "00001101110" => data <= X"AC09639C";
         WHEN "00001101111" => data <= X"00F0A018";
         WHEN "00001110000" => data <= X"00F08018";
         WHEN "00001110001" => data <= X"00F06018";
         WHEN "00001110010" => data <= X"E917A59C";
         WHEN "00001110011" => data <= X"5408849C";
         WHEN "00001110100" => data <= X"1E010000";
         WHEN "00001110101" => data <= X"AC09639C";
         WHEN "00001110110" => data <= X"00F0A018";
         WHEN "00001110111" => data <= X"00F08018";
         WHEN "00001111000" => data <= X"00F06018";
         WHEN "00001111001" => data <= X"EE17A59C";
         WHEN "00001111010" => data <= X"5408849C";
         WHEN "00001111011" => data <= X"17010000";
         WHEN "00001111100" => data <= X"AC09639C";
         WHEN "00001111101" => data <= X"00F0A018";
         WHEN "00001111110" => data <= X"00F08018";
         WHEN "00001111111" => data <= X"00F06018";
         WHEN "00010000000" => data <= X"F317A59C";
         WHEN "00010000001" => data <= X"5408849C";
         WHEN "00010000010" => data <= X"10010000";
         WHEN "00010000011" => data <= X"AC09639C";
         WHEN "00010000100" => data <= X"0000601A";
         WHEN "00010000101" => data <= X"0700A0AA";
         WHEN "00010000110" => data <= X"02A83372";
         WHEN "00010000111" => data <= X"0000E01A";
         WHEN "00010001000" => data <= X"010031A6";
         WHEN "00010001001" => data <= X"00B831E4";
         WHEN "00010001010" => data <= X"FCFFFF13";
         WHEN "00010001011" => data <= X"00000015";
         WHEN "00010001100" => data <= X"00480044";
         WHEN "00010001101" => data <= X"00000015";
         WHEN "00010001110" => data <= X"00006019";
         WHEN "00010001111" => data <= X"02186B71";
         WHEN "00010010000" => data <= X"00480044";
         WHEN "00010010001" => data <= X"00000015";
         WHEN "00010010010" => data <= X"160020AA";
         WHEN "00010010011" => data <= X"02890370";
         WHEN "00010010100" => data <= X"020020AA";
         WHEN "00010010101" => data <= X"070060AA";
         WHEN "00010010110" => data <= X"02991170";
         WHEN "00010010111" => data <= X"EDFFFF03";
         WHEN "00010011000" => data <= X"00000015";
         WHEN "00010011001" => data <= X"E0FF219C";
         WHEN "00010011010" => data <= X"088001D4";
         WHEN "00010011011" => data <= X"0C9001D4";
         WHEN "00010011100" => data <= X"10A001D4";
         WHEN "00010011101" => data <= X"14B001D4";
         WHEN "00010011110" => data <= X"18C001D4";
         WHEN "00010011111" => data <= X"1C4801D4";
         WHEN "00010100000" => data <= X"0000001A";
         WHEN "00010100001" => data <= X"0000401A";
         WHEN "00010100010" => data <= X"160080AA";
         WHEN "00010100011" => data <= X"0100C0AA";
         WHEN "00010100100" => data <= X"070000AB";
         WHEN "00010100101" => data <= X"002092E5";
         WHEN "00010100110" => data <= X"09000010";
         WHEN "00010100111" => data <= X"1C002185";
         WHEN "00010101000" => data <= X"08000186";
         WHEN "00010101001" => data <= X"0C004186";
         WHEN "00010101010" => data <= X"10008186";
         WHEN "00010101011" => data <= X"1400C186";
         WHEN "00010101100" => data <= X"18000187";
         WHEN "00010101101" => data <= X"00480044";
         WHEN "00010101110" => data <= X"2000219C";
         WHEN "00010101111" => data <= X"02A11070";
         WHEN "00010110000" => data <= X"180020AA";
         WHEN "00010110001" => data <= X"008063E2";
         WHEN "00010110010" => data <= X"0000B386";
         WHEN "00010110011" => data <= X"0102B572";
         WHEN "00010110100" => data <= X"02891570";
         WHEN "00010110101" => data <= X"2000A0AA";
         WHEN "00010110110" => data <= X"0100319E";
         WHEN "00010110111" => data <= X"00A831E4";
         WHEN "00010111000" => data <= X"FAFFFF13";
         WHEN "00010111001" => data <= X"0400739E";
         WHEN "00010111010" => data <= X"042001D4";
         WHEN "00010111011" => data <= X"001801D4";
         WHEN "00010111100" => data <= X"02C11670";
         WHEN "00010111101" => data <= X"C7FFFF07";
         WHEN "00010111110" => data <= X"0800529E";
         WHEN "00010111111" => data <= X"2000109E";
         WHEN "00011000000" => data <= X"04008184";
         WHEN "00011000001" => data <= X"E4FFFF03";
         WHEN "00011000010" => data <= X"00006184";
         WHEN "00011000011" => data <= X"B8FF219C";
         WHEN "00011000100" => data <= X"00F08018";
         WHEN "00011000101" => data <= X"2000A0A8";
         WHEN "00011000110" => data <= X"E81E849C";
         WHEN "00011000111" => data <= X"1000619C";
         WHEN "00011001000" => data <= X"308001D4";
         WHEN "00011001001" => data <= X"349001D4";
         WHEN "00011001010" => data <= X"3CB001D4";
         WHEN "00011001011" => data <= X"40C001D4";
         WHEN "00011001100" => data <= X"444801D4";
         WHEN "00011001101" => data <= X"38A001D4";
         WHEN "00011001110" => data <= X"A2010004";
         WHEN "00011001111" => data <= X"00F0401A";
         WHEN "00011010000" => data <= X"00F0001A";
         WHEN "00011010001" => data <= X"5408529E";
         WHEN "00011010010" => data <= X"AC09109E";
         WHEN "00011010011" => data <= X"00F0A018";
         WHEN "00011010100" => data <= X"FC17A59C";
         WHEN "00011010101" => data <= X"049092E0";
         WHEN "00011010110" => data <= X"BC000004";
         WHEN "00011010111" => data <= X"048070E0";
         WHEN "00011011000" => data <= X"1F00201A";
         WHEN "00011011001" => data <= X"00F0A018";
         WHEN "00011011010" => data <= X"0000601A";
         WHEN "00011011011" => data <= X"00FC31AA";
         WHEN "00011011100" => data <= X"0004001B";
         WHEN "00011011101" => data <= X"2000C01A";
         WHEN "00011011110" => data <= X"2D18A59C";
         WHEN "00011011111" => data <= X"0200A0AA";
         WHEN "00011100000" => data <= X"08A891E2";
         WHEN "00011100001" => data <= X"00C094E2";
         WHEN "00011100010" => data <= X"FFFFE0AE";
         WHEN "00011100011" => data <= X"0000B486";
         WHEN "00011100100" => data <= X"00B815E4";
         WHEN "00011100101" => data <= X"1C000010";
         WHEN "00011100110" => data <= X"00000015";
         WHEN "00011100111" => data <= X"0000201A";
         WHEN "00011101000" => data <= X"008813E4";
         WHEN "00011101001" => data <= X"0E000010";
         WHEN "00011101010" => data <= X"049092E0";
         WHEN "00011101011" => data <= X"00F0A018";
         WHEN "00011101100" => data <= X"1F18A59C";
         WHEN "00011101101" => data <= X"049092E0";
         WHEN "00011101110" => data <= X"048070E0";
         WHEN "00011101111" => data <= X"34004186";
         WHEN "00011110000" => data <= X"30000186";
         WHEN "00011110001" => data <= X"38008186";
         WHEN "00011110010" => data <= X"3C00C186";
         WHEN "00011110011" => data <= X"40000187";
         WHEN "00011110100" => data <= X"44002185";
         WHEN "00011110101" => data <= X"9D000000";
         WHEN "00011110110" => data <= X"4800219C";
         WHEN "00011110111" => data <= X"048070E0";
         WHEN "00011111000" => data <= X"9A000004";
         WHEN "00011111001" => data <= X"0C2801D4";
         WHEN "00011111010" => data <= X"98FFFF07";
         WHEN "00011111011" => data <= X"04A074E0";
         WHEN "00011111100" => data <= X"1F00201A";
         WHEN "00011111101" => data <= X"01FC31AA";
         WHEN "00011111110" => data <= X"010060AA";
         WHEN "00011111111" => data <= X"E0FFFF03";
         WHEN "00100000000" => data <= X"0C00A184";
         WHEN "00100000001" => data <= X"0100319E";
         WHEN "00100000010" => data <= X"00B011E4";
         WHEN "00100000011" => data <= X"DDFFFF0F";
         WHEN "00100000100" => data <= X"0200A0AA";
         WHEN "00100000101" => data <= X"00F0A018";
         WHEN "00100000110" => data <= X"4918A59C";
         WHEN "00100000111" => data <= X"049092E0";
         WHEN "00100001000" => data <= X"8A000004";
         WHEN "00100001001" => data <= X"048070E0";
         WHEN "00100001010" => data <= X"1000819E";
         WHEN "00100001011" => data <= X"04A074E2";
         WHEN "00100001100" => data <= X"180020AA";
         WHEN "00100001101" => data <= X"0000B386";
         WHEN "00100001110" => data <= X"0102B572";
         WHEN "00100001111" => data <= X"02891570";
         WHEN "00100010000" => data <= X"2000A0AA";
         WHEN "00100010001" => data <= X"0100319E";
         WHEN "00100010010" => data <= X"00A831E4";
         WHEN "00100010011" => data <= X"FAFFFF13";
         WHEN "00100010100" => data <= X"0400739E";
         WHEN "00100010101" => data <= X"7F00201A";
         WHEN "00100010110" => data <= X"00F031AA";
         WHEN "00100010111" => data <= X"160060AA";
         WHEN "00100011000" => data <= X"02991170";
         WHEN "00100011001" => data <= X"010020AA";
         WHEN "00100011010" => data <= X"070060AA";
         WHEN "00100011011" => data <= X"02991170";
         WHEN "00100011100" => data <= X"68FFFF07";
         WHEN "00100011101" => data <= X"00000015";
         WHEN "00100011110" => data <= X"00F0A018";
         WHEN "00100011111" => data <= X"6A18A59C";
         WHEN "00100100000" => data <= X"049092E0";
         WHEN "00100100001" => data <= X"71000004";
         WHEN "00100100010" => data <= X"048070E0";
         WHEN "00100100011" => data <= X"7F04201A";
         WHEN "00100100100" => data <= X"00F031AA";
         WHEN "00100100101" => data <= X"0000601A";
         WHEN "00100100110" => data <= X"0000B186";
         WHEN "00100100111" => data <= X"0000F486";
         WHEN "00100101000" => data <= X"00A817E4";
         WHEN "00100101001" => data <= X"13000010";
         WHEN "00100101010" => data <= X"0100739E";
         WHEN "00100101011" => data <= X"FFFF739E";
         WHEN "00100101100" => data <= X"00F0A018";
         WHEN "00100101101" => data <= X"08B801D4";
         WHEN "00100101110" => data <= X"04A801D4";
         WHEN "00100101111" => data <= X"009801D4";
         WHEN "00100110000" => data <= X"049092E0";
         WHEN "00100110001" => data <= X"048070E0";
         WHEN "00100110010" => data <= X"60000004";
         WHEN "00100110011" => data <= X"8F18A59C";
         WHEN "00100110100" => data <= X"44002185";
         WHEN "00100110101" => data <= X"30000186";
         WHEN "00100110110" => data <= X"34004186";
         WHEN "00100110111" => data <= X"38008186";
         WHEN "00100111000" => data <= X"3C00C186";
         WHEN "00100111001" => data <= X"40000187";
         WHEN "00100111010" => data <= X"00480044";
         WHEN "00100111011" => data <= X"4800219C";
         WHEN "00100111100" => data <= X"0800A0AA";
         WHEN "00100111101" => data <= X"00A833E4";
         WHEN "00100111110" => data <= X"0400319E";
         WHEN "00100111111" => data <= X"E7FFFF13";
         WHEN "00101000000" => data <= X"0400949E";
         WHEN "00101000001" => data <= X"00F0A018";
         WHEN "00101000010" => data <= X"ABFFFF03";
         WHEN "00101000011" => data <= X"AF18A59C";
         WHEN "00101000100" => data <= X"F0FF219C";
         WHEN "00101000101" => data <= X"048001D4";
         WHEN "00101000110" => data <= X"089001D4";
         WHEN "00101000111" => data <= X"0C4801D4";
         WHEN "00101001000" => data <= X"041843E2";
         WHEN "00101001001" => data <= X"1C0000AA";
         WHEN "00101001010" => data <= X"488024E2";
         WHEN "00101001011" => data <= X"0F0031A6";
         WHEN "00101001100" => data <= X"090060AA";
         WHEN "00101001101" => data <= X"009851E4";
         WHEN "00101001110" => data <= X"03000010";
         WHEN "00101001111" => data <= X"3700719C";
         WHEN "00101010000" => data <= X"3000719C";
         WHEN "00101010001" => data <= X"00900048";
         WHEN "00101010010" => data <= X"002001D4";
         WHEN "00101010011" => data <= X"FCFF109E";
         WHEN "00101010100" => data <= X"FCFF20AE";
         WHEN "00101010101" => data <= X"008830E4";
         WHEN "00101010110" => data <= X"F4FFFF13";
         WHEN "00101010111" => data <= X"00008184";
         WHEN "00101011000" => data <= X"04000186";
         WHEN "00101011001" => data <= X"08004186";
         WHEN "00101011010" => data <= X"0C002185";
         WHEN "00101011011" => data <= X"00480044";
         WHEN "00101011100" => data <= X"1000219C";
         WHEN "00101011101" => data <= X"D4FF219C";
         WHEN "00101011110" => data <= X"0A0020AA";
         WHEN "00101011111" => data <= X"148001D4";
         WHEN "00101100000" => data <= X"189001D4";
         WHEN "00101100001" => data <= X"1CA001D4";
         WHEN "00101100010" => data <= X"24C001D4";
         WHEN "00101100011" => data <= X"041883E2";
         WHEN "00101100100" => data <= X"20B001D4";
         WHEN "00101100101" => data <= X"284801D4";
         WHEN "00101100110" => data <= X"042064E0";
         WHEN "00101100111" => data <= X"0000401A";
         WHEN "00101101000" => data <= X"0000001A";
         WHEN "00101101001" => data <= X"0A00019F";
         WHEN "00101101010" => data <= X"008801D4";
         WHEN "00101101011" => data <= X"041801D4";
         WHEN "00101101100" => data <= X"84040004";
         WHEN "00101101101" => data <= X"00008184";
         WHEN "00101101110" => data <= X"0090D8E2";
         WHEN "00101101111" => data <= X"30006B9D";
         WHEN "00101110000" => data <= X"0000201A";
         WHEN "00101110001" => data <= X"005816D8";
         WHEN "00101110010" => data <= X"008812E4";
         WHEN "00101110011" => data <= X"05000010";
         WHEN "00101110100" => data <= X"04006184";
         WHEN "00101110101" => data <= X"008803E4";
         WHEN "00101110110" => data <= X"04000010";
         WHEN "00101110111" => data <= X"00000015";
         WHEN "00101111000" => data <= X"0100109E";
         WHEN "00101111001" => data <= X"FF0010A6";
         WHEN "00101111010" => data <= X"0100529E";
         WHEN "00101111011" => data <= X"5C040004";
         WHEN "00101111100" => data <= X"00008184";
         WHEN "00101111101" => data <= X"00002186";
         WHEN "00101111110" => data <= X"008832E4";
         WHEN "00101111111" => data <= X"ECFFFF13";
         WHEN "00110000000" => data <= X"04586BE0";
         WHEN "00110000001" => data <= X"0000201A";
         WHEN "00110000010" => data <= X"008830E4";
         WHEN "00110000011" => data <= X"09000010";
         WHEN "00110000100" => data <= X"18004186";
         WHEN "00110000101" => data <= X"14000186";
         WHEN "00110000110" => data <= X"1C008186";
         WHEN "00110000111" => data <= X"2000C186";
         WHEN "00110001000" => data <= X"24000187";
         WHEN "00110001001" => data <= X"28002185";
         WHEN "00110001010" => data <= X"00480044";
         WHEN "00110001011" => data <= X"2C00219C";
         WHEN "00110001100" => data <= X"FFFF109E";
         WHEN "00110001101" => data <= X"008038E2";
         WHEN "00110001110" => data <= X"00A00048";
         WHEN "00110001111" => data <= X"0000718C";
         WHEN "00110010000" => data <= X"F2FFFF03";
         WHEN "00110010001" => data <= X"0000201A";
         WHEN "00110010010" => data <= X"E4FF219C";
         WHEN "00110010011" => data <= X"008001D4";
         WHEN "00110010100" => data <= X"049001D4";
         WHEN "00110010101" => data <= X"08A001D4";
         WHEN "00110010110" => data <= X"0CB001D4";
         WHEN "00110010111" => data <= X"14D001D4";
         WHEN "00110011000" => data <= X"10C001D4";
         WHEN "00110011001" => data <= X"184801D4";
         WHEN "00110011010" => data <= X"041883E2";
         WHEN "00110011011" => data <= X"042004E2";
         WHEN "00110011100" => data <= X"042845E2";
         WHEN "00110011101" => data <= X"1C00C19E";
         WHEN "00110011110" => data <= X"250040AB";
         WHEN "00110011111" => data <= X"00001293";
         WHEN "00110100000" => data <= X"0000201A";
         WHEN "00110100001" => data <= X"008838E4";
         WHEN "00110100010" => data <= X"3C00000C";
         WHEN "00110100011" => data <= X"00D038E4";
         WHEN "00110100100" => data <= X"5B000010";
         WHEN "00110100101" => data <= X"630060AA";
         WHEN "00110100110" => data <= X"01003292";
         WHEN "00110100111" => data <= X"009811E4";
         WHEN "00110101000" => data <= X"4E000010";
         WHEN "00110101001" => data <= X"009851E5";
         WHEN "00110101010" => data <= X"1B000010";
         WHEN "00110101011" => data <= X"0000601A";
         WHEN "00110101100" => data <= X"009811E4";
         WHEN "00110101101" => data <= X"29000010";
         WHEN "00110101110" => data <= X"580060AA";
         WHEN "00110101111" => data <= X"009811E4";
         WHEN "00110110000" => data <= X"37000010";
         WHEN "00110110001" => data <= X"00000015";
         WHEN "00110110010" => data <= X"00A00048";
         WHEN "00110110011" => data <= X"250060A8";
         WHEN "00110110100" => data <= X"0000201A";
         WHEN "00110110101" => data <= X"008810E4";
         WHEN "00110110110" => data <= X"04000010";
         WHEN "00110110111" => data <= X"00000015";
         WHEN "00110111000" => data <= X"00800048";
         WHEN "00110111001" => data <= X"250060A8";
         WHEN "00110111010" => data <= X"0100128F";
         WHEN "00110111011" => data <= X"00A00048";
         WHEN "00110111100" => data <= X"04C078E0";
         WHEN "00110111101" => data <= X"0000201A";
         WHEN "00110111110" => data <= X"008810E4";
         WHEN "00110111111" => data <= X"34000010";
         WHEN "00111000000" => data <= X"00000015";
         WHEN "00111000001" => data <= X"00800048";
         WHEN "00111000010" => data <= X"04C078E0";
         WHEN "00111000011" => data <= X"31000000";
         WHEN "00111000100" => data <= X"0100529E";
         WHEN "00111000101" => data <= X"640060AA";
         WHEN "00111000110" => data <= X"009811E4";
         WHEN "00111000111" => data <= X"EBFFFF0F";
         WHEN "00111001000" => data <= X"00000015";
         WHEN "00111001001" => data <= X"0400169F";
         WHEN "00111001010" => data <= X"04A074E0";
         WHEN "00111001011" => data <= X"0000D686";
         WHEN "00111001100" => data <= X"91FFFF07";
         WHEN "00111001101" => data <= X"04B096E0";
         WHEN "00111001110" => data <= X"0000201A";
         WHEN "00111001111" => data <= X"008810E4";
         WHEN "00111010000" => data <= X"22000010";
         WHEN "00111010001" => data <= X"04B096E0";
         WHEN "00111010010" => data <= X"8BFFFF07";
         WHEN "00111010011" => data <= X"048070E0";
         WHEN "00111010100" => data <= X"1F000000";
         WHEN "00111010101" => data <= X"04C0D8E2";
         WHEN "00111010110" => data <= X"00A00048";
         WHEN "00111010111" => data <= X"04D07AE0";
         WHEN "00111011000" => data <= X"0000201A";
         WHEN "00111011001" => data <= X"008810E4";
         WHEN "00111011010" => data <= X"04000010";
         WHEN "00111011011" => data <= X"04D07AE0";
         WHEN "00111011100" => data <= X"00800048";
         WHEN "00111011101" => data <= X"00000015";
         WHEN "00111011110" => data <= X"00000186";
         WHEN "00111011111" => data <= X"04004186";
         WHEN "00111100000" => data <= X"08008186";
         WHEN "00111100001" => data <= X"0C00C186";
         WHEN "00111100010" => data <= X"10000187";
         WHEN "00111100011" => data <= X"14004187";
         WHEN "00111100100" => data <= X"18002185";
         WHEN "00111100101" => data <= X"00480044";
         WHEN "00111100110" => data <= X"1C00219C";
         WHEN "00111100111" => data <= X"0400169F";
         WHEN "00111101000" => data <= X"04A074E0";
         WHEN "00111101001" => data <= X"0000D686";
         WHEN "00111101010" => data <= X"5AFFFF07";
         WHEN "00111101011" => data <= X"04B096E0";
         WHEN "00111101100" => data <= X"0000201A";
         WHEN "00111101101" => data <= X"008810E4";
         WHEN "00111101110" => data <= X"04000010";
         WHEN "00111101111" => data <= X"04B096E0";
         WHEN "00111110000" => data <= X"54FFFF07";
         WHEN "00111110001" => data <= X"048070E0";
         WHEN "00111110010" => data <= X"04C0D8E2";
         WHEN "00111110011" => data <= X"0100529E";
         WHEN "00111110100" => data <= X"ABFFFF03";
         WHEN "00111110101" => data <= X"0100529E";
         WHEN "00111110110" => data <= X"00005686";
         WHEN "00111110111" => data <= X"00A00048";
         WHEN "00111111000" => data <= X"049072E0";
         WHEN "00111111001" => data <= X"0000201A";
         WHEN "00111111010" => data <= X"008810E4";
         WHEN "00111111011" => data <= X"E3FFFF13";
         WHEN "00111111100" => data <= X"049072E0";
         WHEN "00111111101" => data <= X"DFFFFF03";
         WHEN "00111111110" => data <= X"00000015";
         WHEN "00111111111" => data <= X"00A00048";
         WHEN "01000000000" => data <= X"04C078E0";
         WHEN "01000000001" => data <= X"0000201A";
         WHEN "01000000010" => data <= X"008810E4";
         WHEN "01000000011" => data <= X"F1FFFF13";
         WHEN "01000000100" => data <= X"00000015";
         WHEN "01000000101" => data <= X"00800048";
         WHEN "01000000110" => data <= X"04C078E0";
         WHEN "01000000111" => data <= X"98FFFF03";
         WHEN "01000001000" => data <= X"0100529E";
         WHEN "01000001001" => data <= X"0050201A";
         WHEN "01000001010" => data <= X"030071AA";
         WHEN "01000001011" => data <= X"83FFA0AE";
         WHEN "01000001100" => data <= X"00A813D8";
         WHEN "01000001101" => data <= X"1B00A0AA";
         WHEN "01000001110" => data <= X"00A811D8";
         WHEN "01000001111" => data <= X"010031AA";
         WHEN "01000010000" => data <= X"000011D8";
         WHEN "01000010001" => data <= X"030020AA";
         WHEN "01000010010" => data <= X"008813D8";
         WHEN "01000010011" => data <= X"00480044";
         WHEN "01000010100" => data <= X"00000015";
         WHEN "01000010101" => data <= X"0050601A";
         WHEN "01000010110" => data <= X"0500B3AA";
         WHEN "01000010111" => data <= X"0000358E";
         WHEN "01000011000" => data <= X"400031A6";
         WHEN "01000011001" => data <= X"0000E01A";
         WHEN "01000011010" => data <= X"00B811E4";
         WHEN "01000011011" => data <= X"05000010";
         WHEN "01000011100" => data <= X"00000015";
         WHEN "01000011101" => data <= X"001813D8";
         WHEN "01000011110" => data <= X"00480044";
         WHEN "01000011111" => data <= X"00000015";
         WHEN "01000100000" => data <= X"00000015";
         WHEN "01000100001" => data <= X"F6FFFF03";
         WHEN "01000100010" => data <= X"00000015";
         WHEN "01000100011" => data <= X"0050601A";
         WHEN "01000100100" => data <= X"0500B3AA";
         WHEN "01000100101" => data <= X"0000358E";
         WHEN "01000100110" => data <= X"010031A6";
         WHEN "01000100111" => data <= X"0000E01A";
         WHEN "01000101000" => data <= X"00B811E4";
         WHEN "01000101001" => data <= X"FCFFFF13";
         WHEN "01000101010" => data <= X"00000015";
         WHEN "01000101011" => data <= X"0000738D";
         WHEN "01000101100" => data <= X"00480044";
         WHEN "01000101101" => data <= X"00000015";
         WHEN "01000101110" => data <= X"F8FF219C";
         WHEN "01000101111" => data <= X"FF0063A4";
         WHEN "01000110000" => data <= X"008001D4";
         WHEN "01000110001" => data <= X"D0FF039E";
         WHEN "01000110010" => data <= X"FF0030A6";
         WHEN "01000110011" => data <= X"090060AA";
         WHEN "01000110100" => data <= X"009851E4";
         WHEN "01000110101" => data <= X"0800000C";
         WHEN "01000110110" => data <= X"044801D4";
         WHEN "01000110111" => data <= X"BFFF239E";
         WHEN "01000111000" => data <= X"FF0031A6";
         WHEN "01000111001" => data <= X"050060AA";
         WHEN "01000111010" => data <= X"009851E4";
         WHEN "01000111011" => data <= X"12000010";
         WHEN "01000111100" => data <= X"C9FF039E";
         WHEN "01000111101" => data <= X"E6FFFF07";
         WHEN "01000111110" => data <= X"00000015";
         WHEN "01000111111" => data <= X"FF006BA5";
         WHEN "01001000000" => data <= X"D0FF6B9E";
         WHEN "01001000001" => data <= X"FF00B3A6";
         WHEN "01001000010" => data <= X"0900E0AA";
         WHEN "01001000011" => data <= X"BFFF2B9E";
         WHEN "01001000100" => data <= X"00B855E4";
         WHEN "01001000101" => data <= X"10000010";
         WHEN "01001000110" => data <= X"FF0031A6";
         WHEN "01001000111" => data <= X"040020AA";
         WHEN "01001001000" => data <= X"088810E2";
         WHEN "01001001001" => data <= X"F4FFFF03";
         WHEN "01001001010" => data <= X"008013E2";
         WHEN "01001001011" => data <= X"F2FFFF03";
         WHEN "01001001100" => data <= X"0000001A";
         WHEN "01001001101" => data <= X"9FFF239E";
         WHEN "01001001110" => data <= X"FF0031A6";
         WHEN "01001001111" => data <= X"050060AA";
         WHEN "01001010000" => data <= X"009851E4";
         WHEN "01001010001" => data <= X"FAFFFF13";
         WHEN "01001010010" => data <= X"00000015";
         WHEN "01001010011" => data <= X"EAFFFF03";
         WHEN "01001010100" => data <= X"A9FF039E";
         WHEN "01001010101" => data <= X"050060AA";
         WHEN "01001010110" => data <= X"009851E4";
         WHEN "01001010111" => data <= X"06000010";
         WHEN "01001011000" => data <= X"040020AA";
         WHEN "01001011001" => data <= X"088810E2";
         WHEN "01001011010" => data <= X"C9FF6B9D";
         WHEN "01001011011" => data <= X"E2FFFF03";
         WHEN "01001011100" => data <= X"00800BE2";
         WHEN "01001011101" => data <= X"9FFF2B9E";
         WHEN "01001011110" => data <= X"FF0031A6";
         WHEN "01001011111" => data <= X"050060AA";
         WHEN "01001100000" => data <= X"009851E4";
         WHEN "01001100001" => data <= X"05000010";
         WHEN "01001100010" => data <= X"040020AA";
         WHEN "01001100011" => data <= X"088810E2";
         WHEN "01001100100" => data <= X"F7FFFF03";
         WHEN "01001100101" => data <= X"A9FF6B9D";
         WHEN "01001100110" => data <= X"048070E1";
         WHEN "01001100111" => data <= X"04002185";
         WHEN "01001101000" => data <= X"00000186";
         WHEN "01001101001" => data <= X"00480044";
         WHEN "01001101010" => data <= X"0800219C";
         WHEN "01001101011" => data <= X"FF0063A4";
         WHEN "01001101100" => data <= X"020020AA";
         WHEN "01001101101" => data <= X"00191170";
         WHEN "01001101110" => data <= X"00480044";
         WHEN "01001101111" => data <= X"00000015";
         WHEN "01001110000" => data <= X"041863E1";
         WHEN "01001110001" => data <= X"0000201A";
         WHEN "01001110010" => data <= X"002831E4";
         WHEN "01001110011" => data <= X"04000010";
         WHEN "01001110100" => data <= X"008864E2";
         WHEN "01001110101" => data <= X"00480044";
         WHEN "01001110110" => data <= X"00000015";
         WHEN "01001110111" => data <= X"0000B392";
         WHEN "01001111000" => data <= X"00886BE2";
         WHEN "01001111001" => data <= X"00A813D8";
         WHEN "01001111010" => data <= X"F8FFFF03";
         WHEN "01001111011" => data <= X"0100319E";
         WHEN "01001111100" => data <= X"A8FF219C";
         WHEN "01001111101" => data <= X"00F08018";
         WHEN "01001111110" => data <= X"3800A0A8";
         WHEN "01001111111" => data <= X"081F849C";
         WHEN "01010000000" => data <= X"488001D4";
         WHEN "01010000001" => data <= X"4C9001D4";
         WHEN "01010000010" => data <= X"50A001D4";
         WHEN "01010000011" => data <= X"544801D4";
         WHEN "01010000100" => data <= X"ECFFFF07";
         WHEN "01010000101" => data <= X"1000619C";
         WHEN "01010000110" => data <= X"030020AA";
         WHEN "01010000111" => data <= X"00011170";
         WHEN "01010001000" => data <= X"00F0401A";
         WHEN "01010001001" => data <= X"00F0801A";
         WHEN "01010001010" => data <= X"5408529E";
         WHEN "01010001011" => data <= X"AC09949E";
         WHEN "01010001100" => data <= X"00F0A018";
         WHEN "01010001101" => data <= X"C218A59C";
         WHEN "01010001110" => data <= X"049092E0";
         WHEN "01010001111" => data <= X"03FFFF07";
         WHEN "01010010000" => data <= X"04A074E0";
         WHEN "01010010001" => data <= X"00F0A018";
         WHEN "01010010010" => data <= X"E118A59C";
         WHEN "01010010011" => data <= X"049092E0";
         WHEN "01010010100" => data <= X"FEFEFF07";
         WHEN "01010010101" => data <= X"04A074E0";
         WHEN "01010010110" => data <= X"00F0A018";
         WHEN "01010010111" => data <= X"0419A59C";
         WHEN "01010011000" => data <= X"049092E0";
         WHEN "01010011001" => data <= X"F9FEFF07";
         WHEN "01010011010" => data <= X"04A074E0";
         WHEN "01010011011" => data <= X"FF00201A";
         WHEN "01010011100" => data <= X"FFFF31AA";
         WHEN "01010011101" => data <= X"04000072";
         WHEN "01010011110" => data <= X"0000A01A";
         WHEN "01010011111" => data <= X"038870E2";
         WHEN "01010100000" => data <= X"00A813E4";
         WHEN "01010100001" => data <= X"FCFFFF13";
         WHEN "01010100010" => data <= X"00F0A018";
         WHEN "01010100011" => data <= X"040020AA";
         WHEN "01010100100" => data <= X"488830E2";
         WHEN "01010100101" => data <= X"070031A6";
         WHEN "01010100110" => data <= X"048801D4";
         WHEN "01010100111" => data <= X"070030A6";
         WHEN "01010101000" => data <= X"008801D4";
         WHEN "01010101001" => data <= X"3619A59C";
         WHEN "01010101010" => data <= X"049092E0";
         WHEN "01010101011" => data <= X"E7FEFF07";
         WHEN "01010101100" => data <= X"04A074E0";
         WHEN "01010101101" => data <= X"0C0020AA";
         WHEN "01010101110" => data <= X"488830E2";
         WHEN "01010101111" => data <= X"0F0031A6";
         WHEN "01010110000" => data <= X"0C8801D4";
         WHEN "01010110001" => data <= X"100020AA";
         WHEN "01010110010" => data <= X"488830E2";
         WHEN "01010110011" => data <= X"0F0031A6";
         WHEN "01010110100" => data <= X"088801D4";
         WHEN "01010110101" => data <= X"140020AA";
         WHEN "01010110110" => data <= X"488830E2";
         WHEN "01010110111" => data <= X"0F0031A6";
         WHEN "01010111000" => data <= X"048801D4";
         WHEN "01010111001" => data <= X"180020AA";
         WHEN "01010111010" => data <= X"488830E2";
         WHEN "01010111011" => data <= X"0F0031A6";
         WHEN "01010111100" => data <= X"00F0A018";
         WHEN "01010111101" => data <= X"008801D4";
         WHEN "01010111110" => data <= X"5419A59C";
         WHEN "01010111111" => data <= X"049092E0";
         WHEN "01011000000" => data <= X"D2FEFF07";
         WHEN "01011000001" => data <= X"04A074E0";
         WHEN "01011000010" => data <= X"ADDE201A";
         WHEN "01011000011" => data <= X"0004601A";
         WHEN "01011000100" => data <= X"201431AA";
         WHEN "01011000101" => data <= X"0000B386";
         WHEN "01011000110" => data <= X"008835E4";
         WHEN "01011000111" => data <= X"13000010";
         WHEN "01011001000" => data <= X"0000201A";
         WHEN "01011001001" => data <= X"080010A6";
         WHEN "01011001010" => data <= X"008830E4";
         WHEN "01011001011" => data <= X"0F000010";
         WHEN "01011001100" => data <= X"040033AA";
         WHEN "01011001101" => data <= X"0200A0AA";
         WHEN "01011001110" => data <= X"00003186";
         WHEN "01011001111" => data <= X"08A831E2";
         WHEN "01011010000" => data <= X"008830E4";
         WHEN "01011010001" => data <= X"15000010";
         WHEN "01011010010" => data <= X"0080B3E2";
         WHEN "01011010011" => data <= X"00F0A018";
         WHEN "01011010100" => data <= X"6519A59C";
         WHEN "01011010101" => data <= X"049092E0";
         WHEN "01011010110" => data <= X"BCFEFF07";
         WHEN "01011010111" => data <= X"04A074E0";
         WHEN "01011011000" => data <= X"30000074";
         WHEN "01011011001" => data <= X"00000015";
         WHEN "01011011010" => data <= X"1000019E";
         WHEN "01011011011" => data <= X"0000201A";
         WHEN "01011011100" => data <= X"0000B084";
         WHEN "01011011101" => data <= X"008825E4";
         WHEN "01011011110" => data <= X"0D000010";
         WHEN "01011011111" => data <= X"0400109E";
         WHEN "01011100000" => data <= X"48000186";
         WHEN "01011100001" => data <= X"4C004186";
         WHEN "01011100010" => data <= X"50008186";
         WHEN "01011100011" => data <= X"54002185";
         WHEN "01011100100" => data <= X"00480044";
         WHEN "01011100101" => data <= X"5800219C";
         WHEN "01011100110" => data <= X"0000B586";
         WHEN "01011100111" => data <= X"0400109E";
         WHEN "01011101000" => data <= X"FCAFF0D7";
         WHEN "01011101001" => data <= X"E8FFFF03";
         WHEN "01011101010" => data <= X"008830E4";
         WHEN "01011101011" => data <= X"049092E0";
         WHEN "01011101100" => data <= X"A6FEFF07";
         WHEN "01011101101" => data <= X"04A074E0";
         WHEN "01011101110" => data <= X"EEFFFF03";
         WHEN "01011101111" => data <= X"0000201A";
         WHEN "01011110000" => data <= X"ADDE201A";
         WHEN "01011110001" => data <= X"201471AA";
         WHEN "01011110010" => data <= X"009803E4";
         WHEN "01011110011" => data <= X"14000010";
         WHEN "01011110100" => data <= X"00006019";
         WHEN "01011110101" => data <= X"FFFF601A";
         WHEN "01011110110" => data <= X"039863E0";
         WHEN "01011110111" => data <= X"008823E4";
         WHEN "01011111000" => data <= X"0F000010";
         WHEN "01011111001" => data <= X"FFFF60AD";
         WHEN "01011111010" => data <= X"00F0A018";
         WHEN "01011111011" => data <= X"00F08018";
         WHEN "01011111100" => data <= X"00F06018";
         WHEN "01011111101" => data <= X"FCFF219C";
         WHEN "01011111110" => data <= X"8119A59C";
         WHEN "01011111111" => data <= X"5408849C";
         WHEN "01100000000" => data <= X"004801D4";
         WHEN "01100000001" => data <= X"91FEFF07";
         WHEN "01100000010" => data <= X"AC09639C";
         WHEN "01100000011" => data <= X"FFFF60AD";
         WHEN "01100000100" => data <= X"00002185";
         WHEN "01100000101" => data <= X"00480044";
         WHEN "01100000110" => data <= X"0400219C";
         WHEN "01100000111" => data <= X"00480044";
         WHEN "01100001000" => data <= X"00000015";
         WHEN "01100001001" => data <= X"B0FC219C";
         WHEN "01100001010" => data <= X"247301D4";
         WHEN "01100001011" => data <= X"288301D4";
         WHEN "01100001100" => data <= X"2C9301D4";
         WHEN "01100001101" => data <= X"40E301D4";
         WHEN "01100001110" => data <= X"44F301D4";
         WHEN "01100001111" => data <= X"4C4B01D4";
         WHEN "01100010000" => data <= X"30A301D4";
         WHEN "01100010001" => data <= X"34B301D4";
         WHEN "01100010010" => data <= X"38C301D4";
         WHEN "01100010011" => data <= X"3CD301D4";
         WHEN "01100010100" => data <= X"F5FEFF07";
         WHEN "01100010101" => data <= X"481301D4";
         WHEN "01100010110" => data <= X"66FFFF07";
         WHEN "01100010111" => data <= X"010040AA";
         WHEN "01100011000" => data <= X"00F0201A";
         WHEN "01100011001" => data <= X"701C319E";
         WHEN "01100011010" => data <= X"0000801B";
         WHEN "01100011011" => data <= X"0000C01B";
         WHEN "01100011100" => data <= X"0490D2E1";
         WHEN "01100011101" => data <= X"0000001A";
         WHEN "01100011110" => data <= X"148801D4";
         WHEN "01100011111" => data <= X"04FFFF07";
         WHEN "01100100000" => data <= X"00000015";
         WHEN "01100100001" => data <= X"FF002BA6";
         WHEN "01100100010" => data <= X"270060AA";
         WHEN "01100100011" => data <= X"009811E4";
         WHEN "01100100100" => data <= X"57020010";
         WHEN "01100100101" => data <= X"04580BE3";
         WHEN "01100100110" => data <= X"009851E4";
         WHEN "01100100111" => data <= X"43000010";
         WHEN "01100101000" => data <= X"230060AA";
         WHEN "01100101001" => data <= X"009811E4";
         WHEN "01100101010" => data <= X"82000010";
         WHEN "01100101011" => data <= X"009851E4";
         WHEN "01100101100" => data <= X"10000010";
         WHEN "01100101101" => data <= X"160060AA";
         WHEN "01100101110" => data <= X"F6FF319E";
         WHEN "01100101111" => data <= X"FF0031A6";
         WHEN "01100110000" => data <= X"009851E4";
         WHEN "01100110001" => data <= X"09000010";
         WHEN "01100110010" => data <= X"4000601A";
         WHEN "01100110011" => data <= X"090073AA";
         WHEN "01100110100" => data <= X"488833E2";
         WHEN "01100110101" => data <= X"010031A6";
         WHEN "01100110110" => data <= X"0000601A";
         WHEN "01100110111" => data <= X"009831E4";
         WHEN "01100111000" => data <= X"E7FFFF13";
         WHEN "01100111001" => data <= X"00000015";
         WHEN "01100111010" => data <= X"41000000";
         WHEN "01100111011" => data <= X"00006019";
         WHEN "01100111100" => data <= X"260060AA";
         WHEN "01100111101" => data <= X"009811E4";
         WHEN "01100111110" => data <= X"3D00000C";
         WHEN "01100111111" => data <= X"00006019";
         WHEN "01101000000" => data <= X"E3FEFF07";
         WHEN "01101000001" => data <= X"00004018";
         WHEN "01101000010" => data <= X"00F0A018";
         WHEN "01101000011" => data <= X"00F06018";
         WHEN "01101000100" => data <= X"E319A59C";
         WHEN "01101000101" => data <= X"00008018";
         WHEN "01101000110" => data <= X"AC09639C";
         WHEN "01101000111" => data <= X"4BFEFF07";
         WHEN "01101001000" => data <= X"FF000BA7";
         WHEN "01101001001" => data <= X"200020AA";
         WHEN "01101001010" => data <= X"008818E4";
         WHEN "01101001011" => data <= X"1B000010";
         WHEN "01101001100" => data <= X"2400219E";
         WHEN "01101001101" => data <= X"001042E3";
         WHEN "01101001110" => data <= X"00105AE3";
         WHEN "01101001111" => data <= X"00887AE2";
         WHEN "01101010000" => data <= X"0000201A";
         WHEN "01101010001" => data <= X"0100319E";
         WHEN "01101010010" => data <= X"00C013D8";
         WHEN "01101010011" => data <= X"108801D4";
         WHEN "01101010100" => data <= X"CFFEFF07";
         WHEN "01101010101" => data <= X"0C9801D4";
         WHEN "01101010110" => data <= X"200020AA";
         WHEN "01101010111" => data <= X"FF000BA7";
         WHEN "01101011000" => data <= X"008838E4";
         WHEN "01101011001" => data <= X"0C006186";
         WHEN "01101011010" => data <= X"10002186";
         WHEN "01101011011" => data <= X"F6FFFF13";
         WHEN "01101011100" => data <= X"0100739E";
         WHEN "01101011101" => data <= X"0C037A9E";
         WHEN "01101011110" => data <= X"1800A19E";
         WHEN "01101011111" => data <= X"00A853E3";
         WHEN "01101100000" => data <= X"00885AE3";
         WHEN "01101100001" => data <= X"0100429C";
         WHEN "01101100010" => data <= X"FF0020AA";
         WHEN "01101100011" => data <= X"0088A2E5";
         WHEN "01101100100" => data <= X"BBFFFF0F";
         WHEN "01101100101" => data <= X"0005FADB";
         WHEN "01101100110" => data <= X"BDFEFF07";
         WHEN "01101100111" => data <= X"00000015";
         WHEN "01101101000" => data <= X"E1FFFF03";
         WHEN "01101101001" => data <= X"FF000BA7";
         WHEN "01101101010" => data <= X"2D0060AA";
         WHEN "01101101011" => data <= X"009811E4";
         WHEN "01101101100" => data <= X"0A000010";
         WHEN "01101101101" => data <= X"009851E4";
         WHEN "01101101110" => data <= X"23000010";
         WHEN "01101101111" => data <= X"2A0060AA";
         WHEN "01101110000" => data <= X"009811E4";
         WHEN "01101110001" => data <= X"42000010";
         WHEN "01101110010" => data <= X"2B0060AA";
         WHEN "01101110011" => data <= X"009811E4";
         WHEN "01101110100" => data <= X"0700000C";
         WHEN "01101110101" => data <= X"00006019";
         WHEN "01101110110" => data <= X"ADFEFF07";
         WHEN "01101110111" => data <= X"00000015";
         WHEN "01101111000" => data <= X"180020AA";
         WHEN "01101111001" => data <= X"08886BE1";
         WHEN "01101111010" => data <= X"88886BE1";
         WHEN "01101111011" => data <= X"180060AA";
         WHEN "01101111100" => data <= X"089838E2";
         WHEN "01101111101" => data <= X"889831E2";
         WHEN "01101111110" => data <= X"00004018";
         WHEN "01101111111" => data <= X"2400619E";
         WHEN "01110000000" => data <= X"0000B392";
         WHEN "01110000001" => data <= X"008835E4";
         WHEN "01110000010" => data <= X"06020010";
         WHEN "01110000011" => data <= X"00000015";
         WHEN "01110000100" => data <= X"0100B392";
         WHEN "01110000101" => data <= X"005815E4";
         WHEN "01110000110" => data <= X"0202000C";
         WHEN "01110000111" => data <= X"00F0001B";
         WHEN "01110001000" => data <= X"00F0401B";
         WHEN "01110001001" => data <= X"E11C189F";
         WHEN "01110001010" => data <= X"AC095A9F";
         WHEN "01110001011" => data <= X"0000201A";
         WHEN "01110001100" => data <= X"008832E4";
         WHEN "01110001101" => data <= X"04020010";
         WHEN "01110001110" => data <= X"00000015";
         WHEN "01110001111" => data <= X"90FFFF03";
         WHEN "01110010000" => data <= X"010040AA";
         WHEN "01110010001" => data <= X"3D0060AA";
         WHEN "01110010010" => data <= X"009811E4";
         WHEN "01110010011" => data <= X"E3FFFF13";
         WHEN "01110010100" => data <= X"400060AA";
         WHEN "01110010101" => data <= X"009811E4";
         WHEN "01110010110" => data <= X"E5FFFF0F";
         WHEN "01110010111" => data <= X"00006019";
         WHEN "01110011000" => data <= X"96FEFF07";
         WHEN "01110011001" => data <= X"200060A8";
         WHEN "01110011010" => data <= X"080020AA";
         WHEN "01110011011" => data <= X"00F0A018";
         WHEN "01110011100" => data <= X"00F06018";
         WHEN "01110011101" => data <= X"0888CBE2";
         WHEN "01110011110" => data <= X"005801D4";
         WHEN "01110011111" => data <= X"0A0020AA";
         WHEN "01110100000" => data <= X"F719A59C";
         WHEN "01110100001" => data <= X"00008018";
         WHEN "01110100010" => data <= X"AC09639C";
         WHEN "01110100011" => data <= X"4888D6E2";
         WHEN "01110100100" => data <= X"EEFDFF07";
         WHEN "01110100101" => data <= X"04588BE2";
         WHEN "01110100110" => data <= X"0000201A";
         WHEN "01110100111" => data <= X"008816E4";
         WHEN "01110101000" => data <= X"77FFFF0F";
         WHEN "01110101001" => data <= X"00000015";
         WHEN "01110101010" => data <= X"75FFFF03";
         WHEN "01110101011" => data <= X"0000C01B";
         WHEN "01110101100" => data <= X"00F0A018";
         WHEN "01110101101" => data <= X"D319A59C";
         WHEN "01110101110" => data <= X"00F08018";
         WHEN "01110101111" => data <= X"5408849C";
         WHEN "01110110000" => data <= X"00F06018";
         WHEN "01110110001" => data <= X"25000000";
         WHEN "01110110010" => data <= X"AC09639C";
         WHEN "01110110011" => data <= X"70FEFF07";
         WHEN "01110110100" => data <= X"00000015";
         WHEN "01110110101" => data <= X"FF006BA5";
         WHEN "01110110110" => data <= X"6D0020AA";
         WHEN "01110110111" => data <= X"00880BE4";
         WHEN "01110111000" => data <= X"67010010";
         WHEN "01110111001" => data <= X"00884BE4";
         WHEN "01110111010" => data <= X"39000010";
         WHEN "01110111011" => data <= X"660020AA";
         WHEN "01110111100" => data <= X"00880BE4";
         WHEN "01110111101" => data <= X"E4000010";
         WHEN "01110111110" => data <= X"00884BE4";
         WHEN "01110111111" => data <= X"1B000010";
         WHEN "01111000000" => data <= X"630020AA";
         WHEN "01111000001" => data <= X"00880BE4";
         WHEN "01111000010" => data <= X"9C000010";
         WHEN "01111000011" => data <= X"650020AA";
         WHEN "01111000100" => data <= X"00880BE4";
         WHEN "01111000101" => data <= X"33010010";
         WHEN "01111000110" => data <= X"2A0020AA";
         WHEN "01111000111" => data <= X"00880BE4";
         WHEN "01111001000" => data <= X"57FFFF0F";
         WHEN "01111001001" => data <= X"00000015";
         WHEN "01111001010" => data <= X"00007084";
         WHEN "01111001011" => data <= X"25FFFF07";
         WHEN "01111001100" => data <= X"00000015";
         WHEN "01111001101" => data <= X"0000201A";
         WHEN "01111001110" => data <= X"00F08018";
         WHEN "01111001111" => data <= X"00F06018";
         WHEN "01111010000" => data <= X"00880BE4";
         WHEN "01111010001" => data <= X"5408849C";
         WHEN "01111010010" => data <= X"52000010";
         WHEN "01111010011" => data <= X"AC09639C";
         WHEN "01111010100" => data <= X"00F0A018";
         WHEN "01111010101" => data <= X"151AA59C";
         WHEN "01111010110" => data <= X"BCFDFF07";
         WHEN "01111010111" => data <= X"00000015";
         WHEN "01111011000" => data <= X"47FFFF03";
         WHEN "01111011001" => data <= X"00000015";
         WHEN "01111011010" => data <= X"680020AA";
         WHEN "01111011011" => data <= X"00880BE4";
         WHEN "01111011100" => data <= X"4F000010";
         WHEN "01111011101" => data <= X"690020AA";
         WHEN "01111011110" => data <= X"00880BE4";
         WHEN "01111011111" => data <= X"40FFFF0F";
         WHEN "01111100000" => data <= X"00000015";
         WHEN "01111100001" => data <= X"00007084";
         WHEN "01111100010" => data <= X"0EFFFF07";
         WHEN "01111100011" => data <= X"00000015";
         WHEN "01111100100" => data <= X"0000201A";
         WHEN "01111100101" => data <= X"00880BE4";
         WHEN "01111100110" => data <= X"00F08018";
         WHEN "01111100111" => data <= X"00F06018";
         WHEN "01111101000" => data <= X"04003086";
         WHEN "01111101001" => data <= X"5408849C";
         WHEN "01111101010" => data <= X"58000010";
         WHEN "01111101011" => data <= X"AC09639C";
         WHEN "01111101100" => data <= X"00F0A018";
         WHEN "01111101101" => data <= X"048801D4";
         WHEN "01111101110" => data <= X"000001D4";
         WHEN "01111101111" => data <= X"A3FDFF07";
         WHEN "01111110000" => data <= X"761AA59C";
         WHEN "01111110001" => data <= X"2EFFFF03";
         WHEN "01111110010" => data <= X"00000015";
         WHEN "01111110011" => data <= X"730020AA";
         WHEN "01111110100" => data <= X"00880BE4";
         WHEN "01111110101" => data <= X"40000010";
         WHEN "01111110110" => data <= X"00884BE4";
         WHEN "01111110111" => data <= X"1E000010";
         WHEN "01111111000" => data <= X"700020AA";
         WHEN "01111111001" => data <= X"00880BE4";
         WHEN "01111111010" => data <= X"3F000010";
         WHEN "01111111011" => data <= X"720020AA";
         WHEN "01111111100" => data <= X"00880BE4";
         WHEN "01111111101" => data <= X"22FFFF0F";
         WHEN "01111111110" => data <= X"0004001B";
         WHEN "01111111111" => data <= X"00007884";
         WHEN "10000000000" => data <= X"F0FEFF07";
         WHEN "10000000001" => data <= X"00000015";
         WHEN "10000000010" => data <= X"0000201A";
         WHEN "10000000011" => data <= X"00882BE4";
         WHEN "10000000100" => data <= X"F2000010";
         WHEN "10000000101" => data <= X"00F0A018";
         WHEN "10000000110" => data <= X"040038AA";
         WHEN "10000000111" => data <= X"00007186";
         WHEN "10000001000" => data <= X"020020AA";
         WHEN "10000001001" => data <= X"088873E2";
         WHEN "10000001010" => data <= X"0000201A";
         WHEN "10000001011" => data <= X"009831E4";
         WHEN "10000001100" => data <= X"E5000010";
         WHEN "10000001101" => data <= X"0088B8E2";
         WHEN "10000001110" => data <= X"00F0A018";
         WHEN "10000001111" => data <= X"00F08018";
         WHEN "10000010000" => data <= X"00F06018";
         WHEN "10000010001" => data <= X"6519A59C";
         WHEN "10000010010" => data <= X"5408849C";
         WHEN "10000010011" => data <= X"13000000";
         WHEN "10000010100" => data <= X"AC09639C";
         WHEN "10000010101" => data <= X"740020AA";
         WHEN "10000010110" => data <= X"00880BE4";
         WHEN "10000010111" => data <= X"34000010";
         WHEN "10000011000" => data <= X"760020AA";
         WHEN "10000011001" => data <= X"00880BE4";
         WHEN "10000011010" => data <= X"05FFFF0F";
         WHEN "10000011011" => data <= X"00F0A018";
         WHEN "10000011100" => data <= X"00F08018";
         WHEN "10000011101" => data <= X"00F06018";
         WHEN "10000011110" => data <= X"611AA59C";
         WHEN "10000011111" => data <= X"5408849C";
         WHEN "10000100000" => data <= X"72FDFF07";
         WHEN "10000100001" => data <= X"AC09639C";
         WHEN "10000100010" => data <= X"FDFEFF03";
         WHEN "10000100011" => data <= X"0000C019";
         WHEN "10000100100" => data <= X"00F0A018";
         WHEN "10000100101" => data <= X"301AA59C";
         WHEN "10000100110" => data <= X"6CFDFF07";
         WHEN "10000100111" => data <= X"00000015";
         WHEN "10000101000" => data <= X"30000074";
         WHEN "10000101001" => data <= X"F6FEFF03";
         WHEN "10000101010" => data <= X"00000015";
         WHEN "10000101011" => data <= X"00F0A018";
         WHEN "10000101100" => data <= X"00F06018";
         WHEN "10000101101" => data <= X"311CA59C";
         WHEN "10000101110" => data <= X"00008018";
         WHEN "10000101111" => data <= X"63FDFF07";
         WHEN "10000110000" => data <= X"5408639C";
         WHEN "10000110001" => data <= X"4BFEFF07";
         WHEN "10000110010" => data <= X"00000015";
         WHEN "10000110011" => data <= X"ECFEFF03";
         WHEN "10000110100" => data <= X"00000015";
         WHEN "10000110101" => data <= X"8EFCFF07";
         WHEN "10000110110" => data <= X"00000015";
         WHEN "10000110111" => data <= X"E8FEFF03";
         WHEN "10000111000" => data <= X"00000015";
         WHEN "10000111001" => data <= X"00F0A018";
         WHEN "10000111010" => data <= X"00F08018";
         WHEN "10000111011" => data <= X"00F06018";
         WHEN "10000111100" => data <= X"4D1AA59C";
         WHEN "10000111101" => data <= X"5408849C";
         WHEN "10000111110" => data <= X"54FDFF07";
         WHEN "10000111111" => data <= X"AC09639C";
         WHEN "10001000000" => data <= X"DFFEFF03";
         WHEN "10001000001" => data <= X"0100C0A9";
         WHEN "10001000010" => data <= X"020060AA";
         WHEN "10001000011" => data <= X"089831E2";
         WHEN "10001000100" => data <= X"FFFF319E";
         WHEN "10001000101" => data <= X"00F0A018";
         WHEN "10001000110" => data <= X"008801D4";
         WHEN "10001000111" => data <= X"4BFDFF07";
         WHEN "10001001000" => data <= X"8A1AA59C";
         WHEN "10001001001" => data <= X"D6FEFF03";
         WHEN "10001001010" => data <= X"00000015";
         WHEN "10001001011" => data <= X"0000201A";
         WHEN "10001001100" => data <= X"00F08018";
         WHEN "10001001101" => data <= X"00F06018";
         WHEN "10001001110" => data <= X"008830E4";
         WHEN "10001001111" => data <= X"5408849C";
         WHEN "10001010000" => data <= X"08000010";
         WHEN "10001010001" => data <= X"AC09639C";
         WHEN "10001010010" => data <= X"00F0A018";
         WHEN "10001010011" => data <= X"3FFDFF07";
         WHEN "10001010100" => data <= X"B31AA59C";
         WHEN "10001010101" => data <= X"0000C01B";
         WHEN "10001010110" => data <= X"C9FEFF03";
         WHEN "10001010111" => data <= X"0004001A";
         WHEN "10001011000" => data <= X"00F0A018";
         WHEN "10001011001" => data <= X"39FDFF07";
         WHEN "10001011010" => data <= X"C61AA59C";
         WHEN "10001011011" => data <= X"0000C01B";
         WHEN "10001011100" => data <= X"C3FEFF03";
         WHEN "10001011101" => data <= X"0000001A";
         WHEN "10001011110" => data <= X"0000201A";
         WHEN "10001011111" => data <= X"008810E4";
         WHEN "10001100000" => data <= X"0B000010";
         WHEN "10001100001" => data <= X"00F0A018";
         WHEN "10001100010" => data <= X"00F08018";
         WHEN "10001100011" => data <= X"00F06018";
         WHEN "10001100100" => data <= X"D91AA59C";
         WHEN "10001100101" => data <= X"5408849C";
         WHEN "10001100110" => data <= X"AC09639C";
         WHEN "10001100111" => data <= X"2BFDFF07";
         WHEN "10001101000" => data <= X"0004001A";
         WHEN "10001101001" => data <= X"B6FEFF03";
         WHEN "10001101010" => data <= X"00000015";
         WHEN "10001101011" => data <= X"00007084";
         WHEN "10001101100" => data <= X"84FEFF07";
         WHEN "10001101101" => data <= X"00000015";
         WHEN "10001101110" => data <= X"0000201A";
         WHEN "10001101111" => data <= X"00880BE4";
         WHEN "10001110000" => data <= X"04000010";
         WHEN "10001110001" => data <= X"00F0A018";
         WHEN "10001110010" => data <= X"3CFFFF03";
         WHEN "10001110011" => data <= X"FB1AA59C";
         WHEN "10001110100" => data <= X"3F00201A";
         WHEN "10001110101" => data <= X"FFFF31AA";
         WHEN "10001110110" => data <= X"04007086";
         WHEN "10001110111" => data <= X"0088B3E4";
         WHEN "10001111000" => data <= X"21000010";
         WHEN "10001111001" => data <= X"00F0A018";
         WHEN "10001111010" => data <= X"34FFFF03";
         WHEN "10001111011" => data <= X"181BA59C";
         WHEN "10001111100" => data <= X"0004201A";
         WHEN "10001111101" => data <= X"0088B8E2";
         WHEN "10001111110" => data <= X"00007587";
         WHEN "10001111111" => data <= X"00003887";
         WHEN "10010000000" => data <= X"00C81BE4";
         WHEN "10010000001" => data <= X"10000010";
         WHEN "10010000010" => data <= X"048838E2";
         WHEN "10010000011" => data <= X"00F06018";
         WHEN "10010000100" => data <= X"0000B586";
         WHEN "10010000101" => data <= X"0410A2E0";
         WHEN "10010000110" => data <= X"00003887";
         WHEN "10010000111" => data <= X"04D09AE0";
         WHEN "10010001000" => data <= X"08C801D4";
         WHEN "10010001001" => data <= X"04A801D4";
         WHEN "10010001010" => data <= X"008801D4";
         WHEN "10010001011" => data <= X"AC09639C";
         WHEN "10010001100" => data <= X"10B801D4";
         WHEN "10010001101" => data <= X"05FDFF07";
         WHEN "10010001110" => data <= X"0C9801D4";
         WHEN "10010001111" => data <= X"1000E186";
         WHEN "10010010000" => data <= X"0C006186";
         WHEN "10010010001" => data <= X"0100739E";
         WHEN "10010010010" => data <= X"0400189F";
         WHEN "10010010011" => data <= X"00003786";
         WHEN "10010010100" => data <= X"009851E4";
         WHEN "10010010101" => data <= X"E7FFFF13";
         WHEN "10010010110" => data <= X"00F0A018";
         WHEN "10010010111" => data <= X"17FFFF03";
         WHEN "10010011000" => data <= X"5E1BA59C";
         WHEN "10010011001" => data <= X"00F04018";
         WHEN "10010011010" => data <= X"00F0401B";
         WHEN "10010011011" => data <= X"0000001B";
         WHEN "10010011100" => data <= X"0000601A";
         WHEN "10010011101" => data <= X"0400E0AA";
         WHEN "10010011110" => data <= X"381B429C";
         WHEN "10010011111" => data <= X"F4FFFF03";
         WHEN "10010100000" => data <= X"54085A9F";
         WHEN "10010100001" => data <= X"0000201A";
         WHEN "10010100010" => data <= X"00F0401B";
         WHEN "10010100011" => data <= X"00F0001B";
         WHEN "10010100100" => data <= X"008810E4";
         WHEN "10010100101" => data <= X"54085A9F";
         WHEN "10010100110" => data <= X"07000010";
         WHEN "10010100111" => data <= X"AC09189F";
         WHEN "10010101000" => data <= X"00F0A018";
         WHEN "10010101001" => data <= X"D91AA59C";
         WHEN "10010101010" => data <= X"04D09AE0";
         WHEN "10010101011" => data <= X"BCFFFF03";
         WHEN "10010101100" => data <= X"04C078E0";
         WHEN "10010101101" => data <= X"00007084";
         WHEN "10010101110" => data <= X"42FEFF07";
         WHEN "10010101111" => data <= X"00000015";
         WHEN "10010110000" => data <= X"0000201A";
         WHEN "10010110001" => data <= X"00880BE4";
         WHEN "10010110010" => data <= X"06000010";
         WHEN "10010110011" => data <= X"00F0A018";
         WHEN "10010110100" => data <= X"FB1AA59C";
         WHEN "10010110101" => data <= X"04D09AE0";
         WHEN "10010110110" => data <= X"20FFFF03";
         WHEN "10010110111" => data <= X"04C078E0";
         WHEN "10010111000" => data <= X"3F00201A";
         WHEN "10010111001" => data <= X"FFFF31AA";
         WHEN "10010111010" => data <= X"04007086";
         WHEN "10010111011" => data <= X"0088B3E4";
         WHEN "10010111100" => data <= X"04000010";
         WHEN "10010111101" => data <= X"00F0A018";
         WHEN "10010111110" => data <= X"F7FFFF03";
         WHEN "10010111111" => data <= X"181BA59C";
         WHEN "10011000000" => data <= X"00F0A018";
         WHEN "10011000001" => data <= X"6C1BA59C";
         WHEN "10011000010" => data <= X"04D09AE0";
         WHEN "10011000011" => data <= X"CFFCFF07";
         WHEN "10011000100" => data <= X"04C078E0";
         WHEN "10011000101" => data <= X"00F0A018";
         WHEN "10011000110" => data <= X"0004201A";
         WHEN "10011000111" => data <= X"0000601A";
         WHEN "10011001000" => data <= X"040040A8";
         WHEN "10011001001" => data <= X"00FCE01A";
         WHEN "10011001010" => data <= X"8F1BA59C";
         WHEN "10011001011" => data <= X"0000A286";
         WHEN "10011001100" => data <= X"009855E4";
         WHEN "10011001101" => data <= X"0E000010";
         WHEN "10011001110" => data <= X"FFFF20AF";
         WHEN "10011001111" => data <= X"00F0A018";
         WHEN "10011010000" => data <= X"B61BA59C";
         WHEN "10011010001" => data <= X"04D09AE0";
         WHEN "10011010010" => data <= X"C0FCFF07";
         WHEN "10011010011" => data <= X"04C078E0";
         WHEN "10011010100" => data <= X"00006018";
         WHEN "10011010101" => data <= X"00008284";
         WHEN "10011010110" => data <= X"C3FBFF07";
         WHEN "10011010111" => data <= X"00000015";
         WHEN "10011011000" => data <= X"00F0A018";
         WHEN "10011011001" => data <= X"DCFFFF03";
         WHEN "10011011010" => data <= X"CF1BA59C";
         WHEN "10011011011" => data <= X"0000B186";
         WHEN "10011011100" => data <= X"00C815E4";
         WHEN "10011011101" => data <= X"11000010";
         WHEN "10011011110" => data <= X"00B8B1E2";
         WHEN "10011011111" => data <= X"00A801D4";
         WHEN "10011100000" => data <= X"04D09AE0";
         WHEN "10011100001" => data <= X"04C078E0";
         WHEN "10011100010" => data <= X"209801D4";
         WHEN "10011100011" => data <= X"1CB801D4";
         WHEN "10011100100" => data <= X"188801D4";
         WHEN "10011100101" => data <= X"0C2801D4";
         WHEN "10011100110" => data <= X"ACFCFF07";
         WHEN "10011100111" => data <= X"10A801D4";
         WHEN "10011101000" => data <= X"AAFBFF07";
         WHEN "10011101001" => data <= X"10006184";
         WHEN "10011101010" => data <= X"20006186";
         WHEN "10011101011" => data <= X"1C00E186";
         WHEN "10011101100" => data <= X"18002186";
         WHEN "10011101101" => data <= X"0C00A184";
         WHEN "10011101110" => data <= X"0100739E";
         WHEN "10011101111" => data <= X"DCFFFF03";
         WHEN "10011110000" => data <= X"0400319E";
         WHEN "10011110001" => data <= X"0000B586";
         WHEN "10011110010" => data <= X"0400319E";
         WHEN "10011110011" => data <= X"FCAFF1D7";
         WHEN "10011110100" => data <= X"18FFFF03";
         WHEN "10011110101" => data <= X"009831E4";
         WHEN "10011110110" => data <= X"B8FEFF03";
         WHEN "10011110111" => data <= X"E51BA59C";
         WHEN "10011111000" => data <= X"00F0401B";
         WHEN "10011111001" => data <= X"00F0001B";
         WHEN "10011111010" => data <= X"54085A9F";
         WHEN "10011111011" => data <= X"AC09189F";
         WHEN "10011111100" => data <= X"00F0A018";
         WHEN "10011111101" => data <= X"FB1BA59C";
         WHEN "10011111110" => data <= X"04D09AE0";
         WHEN "10011111111" => data <= X"93FCFF07";
         WHEN "10100000000" => data <= X"04C078E0";
         WHEN "10100000001" => data <= X"00F0A018";
         WHEN "10100000010" => data <= X"00044018";
         WHEN "10100000011" => data <= X"00FCA01A";
         WHEN "10100000100" => data <= X"8F1BA59C";
         WHEN "10100000101" => data <= X"0005601A";
         WHEN "10100000110" => data <= X"FFFFE0AE";
         WHEN "10100000111" => data <= X"00002286";
         WHEN "10100001000" => data <= X"00B811E4";
         WHEN "10100001001" => data <= X"0F000010";
         WHEN "10100001010" => data <= X"00A822E2";
         WHEN "10100001011" => data <= X"008801D4";
         WHEN "10100001100" => data <= X"04D09AE0";
         WHEN "10100001101" => data <= X"04C078E0";
         WHEN "10100001110" => data <= X"1C9801D4";
         WHEN "10100001111" => data <= X"18A801D4";
         WHEN "10100010000" => data <= X"0C2801D4";
         WHEN "10100010001" => data <= X"81FCFF07";
         WHEN "10100010010" => data <= X"108801D4";
         WHEN "10100010011" => data <= X"7FFBFF07";
         WHEN "10100010100" => data <= X"10006184";
         WHEN "10100010101" => data <= X"1C006186";
         WHEN "10100010110" => data <= X"1800A186";
         WHEN "10100010111" => data <= X"0C00A184";
         WHEN "10100011000" => data <= X"0400429C";
         WHEN "10100011001" => data <= X"009822E4";
         WHEN "10100011010" => data <= X"EDFFFF13";
         WHEN "10100011011" => data <= X"FFFFE0AE";
         WHEN "10100011100" => data <= X"00F0A018";
         WHEN "10100011101" => data <= X"98FFFF03";
         WHEN "10100011110" => data <= X"191CA59C";
         WHEN "10100011111" => data <= X"00F0001B";
         WHEN "10100100000" => data <= X"00F0401B";
         WHEN "10100100001" => data <= X"AC09389E";
         WHEN "10100100010" => data <= X"54085A9F";
         WHEN "10100100011" => data <= X"00F0A018";
         WHEN "10100100100" => data <= X"048871E0";
         WHEN "10100100101" => data <= X"341CA59C";
         WHEN "10100100110" => data <= X"04D09AE0";
         WHEN "10100100111" => data <= X"0C8801D4";
         WHEN "10100101000" => data <= X"6AFCFF07";
         WHEN "10100101001" => data <= X"00F0C01B";
         WHEN "10100101010" => data <= X"561C3E9E";
         WHEN "10100101011" => data <= X"0000001B";
         WHEN "10100101100" => data <= X"108801D4";
         WHEN "10100101101" => data <= X"04D09AE0";
         WHEN "10100101110" => data <= X"1000A184";
         WHEN "10100101111" => data <= X"63FCFF07";
         WHEN "10100110000" => data <= X"0C006184";
         WHEN "10100110001" => data <= X"0000201A";
         WHEN "10100110010" => data <= X"0002A01A";
         WHEN "10100110011" => data <= X"020060AA";
         WHEN "10100110100" => data <= X"009818E4";
         WHEN "10100110101" => data <= X"03000010";
         WHEN "10100110110" => data <= X"00000015";
         WHEN "10100110111" => data <= X"0100F172";
         WHEN "10100111000" => data <= X"008811D4";
         WHEN "10100111001" => data <= X"0400319E";
         WHEN "10100111010" => data <= X"00A831E4";
         WHEN "10100111011" => data <= X"F9FFFF13";
         WHEN "10100111100" => data <= X"020060AA";
         WHEN "10100111101" => data <= X"00F0A018";
         WHEN "10100111110" => data <= X"621CA59C";
         WHEN "10100111111" => data <= X"04D09AE0";
         WHEN "10101000000" => data <= X"52FCFF07";
         WHEN "10101000001" => data <= X"0C006184";
         WHEN "10101000010" => data <= X"00004018";
         WHEN "10101000011" => data <= X"0000C01B";
         WHEN "10101000100" => data <= X"0002A01A";
         WHEN "10101000101" => data <= X"020020AA";
         WHEN "10101000110" => data <= X"008818E4";
         WHEN "10101000111" => data <= X"03000010";
         WHEN "10101001000" => data <= X"00000015";
         WHEN "10101001001" => data <= X"0100E272";
         WHEN "10101001010" => data <= X"0000E286";
         WHEN "10101001011" => data <= X"001017E4";
         WHEN "10101001100" => data <= X"12000010";
         WHEN "10101001101" => data <= X"1D0020AA";
         WHEN "10101001110" => data <= X"00885EE4";
         WHEN "10101001111" => data <= X"0E000010";
         WHEN "10101010000" => data <= X"0100FE9E";
         WHEN "10101010001" => data <= X"00002286";
         WHEN "10101010010" => data <= X"04D09AE0";
         WHEN "10101010011" => data <= X"081001D4";
         WHEN "10101010100" => data <= X"048801D4";
         WHEN "10101010101" => data <= X"001001D4";
         WHEN "10101010110" => data <= X"1CA801D4";
         WHEN "10101010111" => data <= X"18B801D4";
         WHEN "10101011000" => data <= X"1400A184";
         WHEN "10101011001" => data <= X"39FCFF07";
         WHEN "10101011010" => data <= X"0C006184";
         WHEN "10101011011" => data <= X"1C00A186";
         WHEN "10101011100" => data <= X"1800E186";
         WHEN "10101011101" => data <= X"04B8D7E3";
         WHEN "10101011110" => data <= X"0400429C";
         WHEN "10101011111" => data <= X"00A822E4";
         WHEN "10101100000" => data <= X"E6FFFF13";
         WHEN "10101100001" => data <= X"020020AA";
         WHEN "10101100010" => data <= X"0000201A";
         WHEN "10101100011" => data <= X"00881EE4";
         WHEN "10101100100" => data <= X"11000010";
         WHEN "10101100101" => data <= X"0100189F";
         WHEN "10101100110" => data <= X"FFFF189F";
         WHEN "10101100111" => data <= X"00F0A018";
         WHEN "10101101000" => data <= X"00F001D4";
         WHEN "10101101001" => data <= X"8C1CA59C";
         WHEN "10101101010" => data <= X"04D09AE0";
         WHEN "10101101011" => data <= X"27FCFF07";
         WHEN "10101101100" => data <= X"0C006184";
         WHEN "10101101101" => data <= X"00F0A018";
         WHEN "10101101110" => data <= X"00F001D4";
         WHEN "10101101111" => data <= X"A51CA59C";
         WHEN "10101110000" => data <= X"04D09AE0";
         WHEN "10101110001" => data <= X"21FCFF07";
         WHEN "10101110010" => data <= X"0C006184";
         WHEN "10101110011" => data <= X"ACFDFF03";
         WHEN "10101110100" => data <= X"0000C01B";
         WHEN "10101110101" => data <= X"030020AA";
         WHEN "10101110110" => data <= X"008838E4";
         WHEN "10101110111" => data <= X"B7FFFF13";
         WHEN "10101111000" => data <= X"04D09AE0";
         WHEN "10101111001" => data <= X"F5FFFF03";
         WHEN "10101111010" => data <= X"00F0A018";
         WHEN "10101111011" => data <= X"A8FCFF07";
         WHEN "10101111100" => data <= X"00000015";
         WHEN "10101111101" => data <= X"A6FCFF07";
         WHEN "10101111110" => data <= X"FF000BA7";
         WHEN "10101111111" => data <= X"D0FF189F";
         WHEN "10110000000" => data <= X"020020AA";
         WHEN "10110000001" => data <= X"088838E2";
         WHEN "10110000010" => data <= X"FF004BA6";
         WHEN "10110000011" => data <= X"00C031E2";
         WHEN "10110000100" => data <= X"008831E2";
         WHEN "10110000101" => data <= X"D0FF529E";
         WHEN "10110000110" => data <= X"99FDFF03";
         WHEN "10110000111" => data <= X"008852E2";
         WHEN "10110001000" => data <= X"0100429C";
         WHEN "10110001001" => data <= X"0001A0AA";
         WHEN "10110001010" => data <= X"00A822E4";
         WHEN "10110001011" => data <= X"F5FDFF13";
         WHEN "10110001100" => data <= X"0300739E";
         WHEN "10110001101" => data <= X"00F0A018";
         WHEN "10110001110" => data <= X"1F1DA59C";
         WHEN "10110001111" => data <= X"21FEFF03";
         WHEN "10110010000" => data <= X"00008018";
         WHEN "10110010001" => data <= X"00881CE4";
         WHEN "10110010010" => data <= X"18000010";
         WHEN "10110010011" => data <= X"080020AA";
         WHEN "10110010100" => data <= X"088894E2";
         WHEN "10110010101" => data <= X"01009C9F";
         WHEN "10110010110" => data <= X"040020AA";
         WHEN "10110010111" => data <= X"00883CE4";
         WHEN "10110011000" => data <= X"2E000010";
         WHEN "10110011001" => data <= X"00A082E2";
         WHEN "10110011010" => data <= X"0000201A";
         WHEN "10110011011" => data <= X"008810E4";
         WHEN "10110011100" => data <= X"10000010";
         WHEN "10110011101" => data <= X"0000601A";
         WHEN "10110011110" => data <= X"008836E4";
         WHEN "10110011111" => data <= X"80FDFF13";
         WHEN "10110100000" => data <= X"010040AA";
         WHEN "10110100001" => data <= X"00F0A018";
         WHEN "10110100010" => data <= X"00F08018";
         WHEN "10110100011" => data <= X"00F06018";
         WHEN "10110100100" => data <= X"C01CA59C";
         WHEN "10110100101" => data <= X"5408849C";
         WHEN "10110100110" => data <= X"ECFBFF07";
         WHEN "10110100111" => data <= X"AC09639C";
         WHEN "10110101000" => data <= X"77FDFF03";
         WHEN "10110101001" => data <= X"0490D2E2";
         WHEN "10110101010" => data <= X"EBFFFF03";
         WHEN "10110101011" => data <= X"0000801A";
         WHEN "10110101100" => data <= X"020020AA";
         WHEN "10110101101" => data <= X"088896E3";
         WHEN "10110101110" => data <= X"FF3F36A6";
         WHEN "10110101111" => data <= X"009831E4";
         WHEN "10110110000" => data <= X"06000010";
         WHEN "10110110001" => data <= X"04C0B8E0";
         WHEN "10110110010" => data <= X"00E001D4";
         WHEN "10110110011" => data <= X"00008018";
         WHEN "10110110100" => data <= X"DEFBFF07";
         WHEN "10110110101" => data <= X"04D07AE0";
         WHEN "10110110110" => data <= X"0000201A";
         WHEN "10110110111" => data <= X"00880EE4";
         WHEN "10110111000" => data <= X"10000010";
         WHEN "10110111001" => data <= X"00E030E2";
         WHEN "10110111010" => data <= X"01007472";
         WHEN "10110111011" => data <= X"009811D4";
         WHEN "10110111100" => data <= X"0100D69E";
         WHEN "10110111101" => data <= X"00B07EE4";
         WHEN "10110111110" => data <= X"07000010";
         WHEN "10110111111" => data <= X"0000201A";
         WHEN "10111000000" => data <= X"00880EE4";
         WHEN "10111000001" => data <= X"04000010";
         WHEN "10111000010" => data <= X"00000015";
         WHEN "10111000011" => data <= X"04B010D4";
         WHEN "10111000100" => data <= X"04B0D6E3";
         WHEN "10111000101" => data <= X"0000801B";
         WHEN "10111000110" => data <= X"C5FDFF03";
         WHEN "10111000111" => data <= X"FFFF529E";
         WHEN "10111001000" => data <= X"00003186";
         WHEN "10111001001" => data <= X"01003172";
         WHEN "10111001010" => data <= X"008814E4";
         WHEN "10111001011" => data <= X"F1FFFF13";
         WHEN "10111001100" => data <= X"00F0A018";
         WHEN "10111001101" => data <= X"00F06018";
         WHEN "10111001110" => data <= X"08A001D4";
         WHEN "10111001111" => data <= X"048801D4";
         WHEN "10111010000" => data <= X"00E001D4";
         WHEN "10111010001" => data <= X"F41CA59C";
         WHEN "10111010010" => data <= X"00008018";
         WHEN "10111010011" => data <= X"BFFBFF07";
         WHEN "10111010100" => data <= X"AC09639C";
         WHEN "10111010101" => data <= X"E8FFFF03";
         WHEN "10111010110" => data <= X"0100D69E";
         WHEN "10111010111" => data <= X"000004E4";
         WHEN "10111011000" => data <= X"000060A9";
         WHEN "10111011001" => data <= X"15000010";
         WHEN "10111011010" => data <= X"000083A9";
         WHEN "10111011011" => data <= X"0100C0A8";
         WHEN "10111011100" => data <= X"000084E5";
         WHEN "10111011101" => data <= X"05000010";
         WHEN "10111011110" => data <= X"006084E4";
         WHEN "10111011111" => data <= X"002084E0";
         WHEN "10111100000" => data <= X"FCFFFF13";
         WHEN "10111100001" => data <= X"0030C6E0";
         WHEN "10111100010" => data <= X"0030EBE0";
         WHEN "10111100011" => data <= X"4100C6B8";
         WHEN "10111100100" => data <= X"02200CE1";
         WHEN "10111100101" => data <= X"0060A4E4";
         WHEN "10111100110" => data <= X"410084B8";
         WHEN "10111100111" => data <= X"0400000C";
         WHEN "10111101000" => data <= X"00000015";
         WHEN "10111101001" => data <= X"000067A9";
         WHEN "10111101010" => data <= X"000088A9";
         WHEN "10111101011" => data <= X"000026E4";
         WHEN "10111101100" => data <= X"F7FFFF13";
         WHEN "10111101101" => data <= X"0030EBE0";
         WHEN "10111101110" => data <= X"00480044";
         WHEN "10111101111" => data <= X"00000015";
         WHEN "10111110000" => data <= X"0000A9A9";
         WHEN "10111110001" => data <= X"E6FFFF07";
         WHEN "10111110010" => data <= X"00000015";
         WHEN "10111110011" => data <= X"00680044";
         WHEN "10111110100" => data <= X"00006CA9";
         WHEN "10111110101" => data <= X"65202449";
         WHEN "10111110110" => data <= X"726F7272";
         WHEN "10111110111" => data <= X"44000A21";
         WHEN "10111111000" => data <= X"72652024";
         WHEN "10111111001" => data <= X"0A726F72";
         WHEN "10111111010" => data <= X"71726900";
         WHEN "10111111011" => data <= X"3F3F000A";
         WHEN "10111111100" => data <= X"73000A3F";
         WHEN "10111111101" => data <= X"65747379";
         WHEN "10111111110" => data <= X"000A216D";
         WHEN "10111111111" => data <= X"63656843";
         WHEN "11000000000" => data <= X"676E696B";
         WHEN "11000000001" => data <= X"73616C20";
         WHEN "11000000010" => data <= X"61702074";
         WHEN "11000000011" => data <= X"6F206567";
         WHEN "11000000100" => data <= X"6C662066";
         WHEN "11000000101" => data <= X"20687361";
         WHEN "11000000110" => data <= X"74706D65";
         WHEN "11000000111" => data <= X"46000A79";
         WHEN "11000001000" => data <= X"6873616C";
         WHEN "11000001001" => data <= X"72726520";
         WHEN "11000001010" => data <= X"0A21726F";
         WHEN "11000001011" => data <= X"61724500";
         WHEN "11000001100" => data <= X"676E6973";
         WHEN "11000001101" => data <= X"73616C20";
         WHEN "11000001110" => data <= X"61702074";
         WHEN "11000001111" => data <= X"6F206567";
         WHEN "11000010000" => data <= X"6C462066";
         WHEN "11000010001" => data <= X"0A687361";
         WHEN "11000010010" => data <= X"69725700";
         WHEN "11000010011" => data <= X"676E6974";
         WHEN "11000010100" => data <= X"73657420";
         WHEN "11000010101" => data <= X"65732074";
         WHEN "11000010110" => data <= X"6E657571";
         WHEN "11000010111" => data <= X"74206563";
         WHEN "11000011000" => data <= X"6C66206F";
         WHEN "11000011001" => data <= X"2E687361";
         WHEN "11000011010" => data <= X"6556000A";
         WHEN "11000011011" => data <= X"79666972";
         WHEN "11000011100" => data <= X"20676E69";
         WHEN "11000011101" => data <= X"74736574";
         WHEN "11000011110" => data <= X"71657320";
         WHEN "11000011111" => data <= X"636E6575";
         WHEN "11000100000" => data <= X"72662065";
         WHEN "11000100001" => data <= X"66206D6F";
         WHEN "11000100010" => data <= X"6873616C";
         WHEN "11000100011" => data <= X"54000A2E";
         WHEN "11000100100" => data <= X"20747365";
         WHEN "11000100101" => data <= X"6C696166";
         WHEN "11000100110" => data <= X"203A6465";
         WHEN "11000100111" => data <= X"3A206425";
         WHEN "11000101000" => data <= X"25783020";
         WHEN "11000101001" => data <= X"3D2F2058";
         WHEN "11000101010" => data <= X"25783020";
         WHEN "11000101011" => data <= X"46000A58";
         WHEN "11000101100" => data <= X"6873616C";
         WHEN "11000101101" => data <= X"73657420";
         WHEN "11000101110" => data <= X"6B6F2074";
         WHEN "11000101111" => data <= X"0A2E7961";
         WHEN "11000110000" => data <= X"5343000A";
         WHEN "11000110001" => data <= X"3637342D";
         WHEN "11000110010" => data <= X"626D4520";
         WHEN "11000110011" => data <= X"65646465";
         WHEN "11000110100" => data <= X"79532064";
         WHEN "11000110101" => data <= X"6D657473";
         WHEN "11000110110" => data <= X"73654420";
         WHEN "11000110111" => data <= X"0A6E6769";
         WHEN "11000111000" => data <= X"65704F00";
         WHEN "11000111001" => data <= X"7369726E";
         WHEN "11000111010" => data <= X"61622063";
         WHEN "11000111011" => data <= X"20646573";
         WHEN "11000111100" => data <= X"74726976";
         WHEN "11000111101" => data <= X"206C6175";
         WHEN "11000111110" => data <= X"746F7250";
         WHEN "11000111111" => data <= X"7079746F";
         WHEN "11001000000" => data <= X"000A2E65";
         WHEN "11001000001" => data <= X"6C697542";
         WHEN "11001000010" => data <= X"65762064";
         WHEN "11001000011" => data <= X"6F697372";
         WHEN "11001000100" => data <= X"53203A6E";
         WHEN "11001000101" => data <= X"41206E75";
         WHEN "11001000110" => data <= X"31206775";
         WHEN "11001000111" => data <= X"30312030";
         WHEN "11001001000" => data <= X"3A36353A";
         WHEN "11001001001" => data <= X"41203130";
         WHEN "11001001010" => data <= X"4543204D";
         WHEN "11001001011" => data <= X"32205453";
         WHEN "11001001100" => data <= X"0A353230";
         WHEN "11001001101" => data <= X"2049000A";
         WHEN "11001001110" => data <= X"43206D61";
         WHEN "11001001111" => data <= X"25205550";
         WHEN "11001010000" => data <= X"666F2064";
         WHEN "11001010001" => data <= X"20642520";
         WHEN "11001010010" => data <= X"6E6E7572";
         WHEN "11001010011" => data <= X"20676E69";
         WHEN "11001010100" => data <= X"00207461";
         WHEN "11001010101" => data <= X"64256425";
         WHEN "11001010110" => data <= X"2564252E";
         WHEN "11001010111" => data <= X"484D2064";
         WHEN "11001011000" => data <= X"0A0A2E7A";
         WHEN "11001011001" => data <= X"65784500";
         WHEN "11001011010" => data <= X"69747563";
         WHEN "11001011011" => data <= X"6620676E";
         WHEN "11001011100" => data <= X"6873616C";
         WHEN "11001011101" => data <= X"6F727020";
         WHEN "11001011110" => data <= X"6D617267";
         WHEN "11001011111" => data <= X"0A2E2E2E";
         WHEN "11001100000" => data <= X"6F725000";
         WHEN "11001100001" => data <= X"6D617267";
         WHEN "11001100010" => data <= X"65727020";
         WHEN "11001100011" => data <= X"746E6573";
         WHEN "11001100100" => data <= X"74756220";
         WHEN "11001100101" => data <= X"746F6E20";
         WHEN "11001100110" => data <= X"726F6620";
         WHEN "11001100111" => data <= X"69687420";
         WHEN "11001101000" => data <= X"61542073";
         WHEN "11001101001" => data <= X"74656772";
         WHEN "11001101010" => data <= X"69440A2E";
         WHEN "11001101011" => data <= X"6F792064";
         WHEN "11001101100" => data <= X"70752075";
         WHEN "11001101101" => data <= X"64616F6C";
         WHEN "11001101110" => data <= X"726F6620";
         WHEN "11001101111" => data <= X"65687420";
         WHEN "11001110000" => data <= X"31524F20";
         WHEN "11001110001" => data <= X"20303234";
         WHEN "11001110010" => data <= X"74616C70";
         WHEN "11001110011" => data <= X"6D726F66";
         WHEN "11001110100" => data <= X"44000A3F";
         WHEN "11001110101" => data <= X"6C6E776F";
         WHEN "11001110110" => data <= X"3A64616F";
         WHEN "11001110111" => data <= X"6E6F6420";
         WHEN "11001111000" => data <= X"52000A65";
         WHEN "11001111001" => data <= X"69646165";
         WHEN "11001111010" => data <= X"6320676E";
         WHEN "11001111011" => data <= X"2065646F";
         WHEN "11001111100" => data <= X"6C626174";
         WHEN "11001111101" => data <= X"44000A65";
         WHEN "11001111110" => data <= X"6C6E776F";
         WHEN "11001111111" => data <= X"3A64616F";
         WHEN "11010000000" => data <= X"74657320";
         WHEN "11010000001" => data <= X"64646120";
         WHEN "11010000010" => data <= X"73736572";
         WHEN "11010000011" => data <= X"30203D20";
         WHEN "11010000100" => data <= X"0A582578";
         WHEN "11010000101" => data <= X"72724500";
         WHEN "11010000110" => data <= X"202C726F";
         WHEN "11010000111" => data <= X"70206F6E";
         WHEN "11010001000" => data <= X"72676F72";
         WHEN "11010001001" => data <= X"6C206D61";
         WHEN "11010001010" => data <= X"6564616F";
         WHEN "11010001011" => data <= X"000A2164";
         WHEN "11010001100" => data <= X"63657845";
         WHEN "11010001101" => data <= X"6E697475";
         WHEN "11010001110" => data <= X"6F6C2067";
         WHEN "11010001111" => data <= X"64656461";
         WHEN "11010010000" => data <= X"6F727020";
         WHEN "11010010001" => data <= X"6D617267";
         WHEN "11010010010" => data <= X"0A2E2E2E";
         WHEN "11010010011" => data <= X"74655300";
         WHEN "11010010100" => data <= X"676E6974";
         WHEN "11010010101" => data <= X"6F727020";
         WHEN "11010010110" => data <= X"6D202E67";
         WHEN "11010010111" => data <= X"0A65646F";
         WHEN "11010011000" => data <= X"74655300";
         WHEN "11010011001" => data <= X"676E6974";
         WHEN "11010011010" => data <= X"72657620";
         WHEN "11010011011" => data <= X"202E6669";
         WHEN "11010011100" => data <= X"65646F6D";
         WHEN "11010011101" => data <= X"6F4E000A";
         WHEN "11010011110" => data <= X"6F727020";
         WHEN "11010011111" => data <= X"6D617267";
         WHEN "11010100000" => data <= X"65727020";
         WHEN "11010100001" => data <= X"746E6573";
         WHEN "11010100010" => data <= X"7250000A";
         WHEN "11010100011" => data <= X"6172676F";
         WHEN "11010100100" => data <= X"6E69206D";
         WHEN "11010100101" => data <= X"6D656D20";
         WHEN "11010100110" => data <= X"6F726620";
         WHEN "11010100111" => data <= X"6162206D";
         WHEN "11010101000" => data <= X"302B6573";
         WHEN "11010101001" => data <= X"206F7420";
         WHEN "11010101010" => data <= X"65736162";
         WHEN "11010101011" => data <= X"2578302B";
         WHEN "11010101100" => data <= X"53000A58";
         WHEN "11010101101" => data <= X"63746977";
         WHEN "11010101110" => data <= X"20646568";
         WHEN "11010101111" => data <= X"46206F74";
         WHEN "11010110000" => data <= X"6873616C";
         WHEN "11010110001" => data <= X"7753000A";
         WHEN "11010110010" => data <= X"68637469";
         WHEN "11010110011" => data <= X"74206465";
         WHEN "11010110100" => data <= X"4453206F";
         WHEN "11010110101" => data <= X"0A6D6152";
         WHEN "11010110110" => data <= X"656C5000";
         WHEN "11010110111" => data <= X"20657361";
         WHEN "11010111000" => data <= X"6E616863";
         WHEN "11010111001" => data <= X"74206567";
         WHEN "11010111010" => data <= X"6874206F";
         WHEN "11010111011" => data <= X"44532065";
         WHEN "11010111100" => data <= X"204D4152";
         WHEN "11010111101" => data <= X"2A207962";
         WHEN "11010111110" => data <= X"4E000A74";
         WHEN "11010111111" => data <= X"7270206F";
         WHEN "11011000000" => data <= X"6172676F";
         WHEN "11011000001" => data <= X"6F6C206D";
         WHEN "11011000010" => data <= X"64656461";
         WHEN "11011000011" => data <= X"206E6920";
         WHEN "11011000100" => data <= X"61524453";
         WHEN "11011000101" => data <= X"000A216D";
         WHEN "11011000110" => data <= X"676F7250";
         WHEN "11011000111" => data <= X"206D6172";
         WHEN "11011001000" => data <= X"73656F64";
         WHEN "11011001001" => data <= X"746F6E20";
         WHEN "11011001010" => data <= X"74696620";
         WHEN "11011001011" => data <= X"206E6920";
         WHEN "11011001100" => data <= X"73616C46";
         WHEN "11011001101" => data <= X"000A2168";
         WHEN "11011001110" => data <= X"706D6F43";
         WHEN "11011001111" => data <= X"20657261";
         WHEN "11011010000" => data <= X"6F727265";
         WHEN "11011010001" => data <= X"74612072";
         WHEN "11011010010" => data <= X"25783020";
         WHEN "11011010011" => data <= X"203A2058";
         WHEN "11011010100" => data <= X"58257830";
         WHEN "11011010101" => data <= X"203D2120";
         WHEN "11011010110" => data <= X"58257830";
         WHEN "11011010111" => data <= X"6F43000A";
         WHEN "11011011000" => data <= X"7261706D";
         WHEN "11011011001" => data <= X"6F642065";
         WHEN "11011011010" => data <= X"000A656E";
         WHEN "11011011011" => data <= X"63656843";
         WHEN "11011011100" => data <= X"676E696B";
         WHEN "11011011101" => data <= X"20666920";
         WHEN "11011011110" => data <= X"20656874";
         WHEN "11011011111" => data <= X"73616C66";
         WHEN "11011100000" => data <= X"73692068";
         WHEN "11011100001" => data <= X"706D6520";
         WHEN "11011100010" => data <= X"2E2E7974";
         WHEN "11011100011" => data <= X"53000A2E";
         WHEN "11011100100" => data <= X"74726174";
         WHEN "11011100101" => data <= X"616C6620";
         WHEN "11011100110" => data <= X"65206873";
         WHEN "11011100111" => data <= X"65736172";
         WHEN "11011101000" => data <= X"63796320";
         WHEN "11011101001" => data <= X"6620656C";
         WHEN "11011101010" => data <= X"7020726F";
         WHEN "11011101011" => data <= X"20656761";
         WHEN "11011101100" => data <= X"58257830";
         WHEN "11011101101" => data <= X"7453000A";
         WHEN "11011101110" => data <= X"20747261";
         WHEN "11011101111" => data <= X"676F7270";
         WHEN "11011110000" => data <= X"6D6D6172";
         WHEN "11011110001" => data <= X"20676E69";
         WHEN "11011110010" => data <= X"73616C66";
         WHEN "11011110011" => data <= X"50000A68";
         WHEN "11011110100" => data <= X"72676F72";
         WHEN "11011110101" => data <= X"696D6D61";
         WHEN "11011110110" => data <= X"6620676E";
         WHEN "11011110111" => data <= X"73696E69";
         WHEN "11011111000" => data <= X"0A646568";
         WHEN "11011111001" => data <= X"206F4E00";
         WHEN "11011111010" => data <= X"676F7270";
         WHEN "11011111011" => data <= X"206D6172";
         WHEN "11011111100" => data <= X"66206E69";
         WHEN "11011111101" => data <= X"6873616C";
         WHEN "11011111110" => data <= X"43000A21";
         WHEN "11011111111" => data <= X"6B636568";
         WHEN "11100000000" => data <= X"20676E69";
         WHEN "11100000001" => data <= X"66206669";
         WHEN "11100000010" => data <= X"6873616C";
         WHEN "11100000011" => data <= X"20736920";
         WHEN "11100000100" => data <= X"72696427";
         WHEN "11100000101" => data <= X"0A277974";
         WHEN "11100000110" => data <= X"616C4600";
         WHEN "11100000111" => data <= X"69206873";
         WHEN "11100001000" => data <= X"6D652073";
         WHEN "11100001001" => data <= X"20797470";
         WHEN "11100001010" => data <= X"61726528";
         WHEN "11100001011" => data <= X"29646573";
         WHEN "11100001100" => data <= X"000A0A2E";
         WHEN "11100001101" => data <= X"72617453";
         WHEN "11100001110" => data <= X"676E6974";
         WHEN "11100001111" => data <= X"6D697320";
         WHEN "11100010000" => data <= X"20656C70";
         WHEN "11100010001" => data <= X"61524453";
         WHEN "11100010010" => data <= X"656D206D";
         WHEN "11100010011" => data <= X"6568636D";
         WHEN "11100010100" => data <= X"0A2E6B63";
         WHEN "11100010101" => data <= X"7257000A";
         WHEN "11100010110" => data <= X"6E697469";
         WHEN "11100010111" => data <= X"2E2E2E67";
         WHEN "11100011000" => data <= X"6556000A";
         WHEN "11100011001" => data <= X"79666972";
         WHEN "11100011010" => data <= X"2E676E69";
         WHEN "11100011011" => data <= X"000A2E2E";
         WHEN "11100011100" => data <= X"6F727245";
         WHEN "11100011101" => data <= X"30402072";
         WHEN "11100011110" => data <= X"20582578";
         WHEN "11100011111" => data <= X"7830203A";
         WHEN "11100100000" => data <= X"21205825";
         WHEN "11100100001" => data <= X"7830203D";
         WHEN "11100100010" => data <= X"000A5825";
         WHEN "11100100011" => data <= X"6F20724E";
         WHEN "11100100100" => data <= X"72652066";
         WHEN "11100100101" => data <= X"73726F72";
         WHEN "11100100110" => data <= X"756F6620";
         WHEN "11100100111" => data <= X"3A20646E";
         WHEN "11100101000" => data <= X"0A642520";
         WHEN "11100101001" => data <= X"6D654D00";
         WHEN "11100101010" => data <= X"63656863";
         WHEN "11100101011" => data <= X"6F64206B";
         WHEN "11100101100" => data <= X"202C656E";
         WHEN "11100101101" => data <= X"65206425";
         WHEN "11100101110" => data <= X"726F7272";
         WHEN "11100101111" => data <= X"000A0A73";
         WHEN "11100110000" => data <= X"6E6E6143";
         WHEN "11100110001" => data <= X"7020746F";
         WHEN "11100110010" => data <= X"72676F72";
         WHEN "11100110011" => data <= X"66206D61";
         WHEN "11100110100" => data <= X"6873616C";
         WHEN "11100110101" => data <= X"6261202C";
         WHEN "11100110110" => data <= X"6974726F";
         WHEN "11100110111" => data <= X"0A21676E";
         WHEN "11100111000" => data <= X"776F4400";
         WHEN "11100111001" => data <= X"616F6C6E";
         WHEN "11100111010" => data <= X"61203A64";
         WHEN "11100111011" => data <= X"78302074";
         WHEN "11100111100" => data <= X"000A5825";
         WHEN "11100111101" => data <= X"69726556";
         WHEN "11100111110" => data <= X"61636966";
         WHEN "11100111111" => data <= X"6E6F6974";
         WHEN "11101000000" => data <= X"72726520";
         WHEN "11101000001" => data <= X"6120726F";
         WHEN "11101000010" => data <= X"78302074";
         WHEN "11101000011" => data <= X"3A205825";
         WHEN "11101000100" => data <= X"25783020";
         WHEN "11101000101" => data <= X"3D212058";
         WHEN "11101000110" => data <= X"25783020";
         WHEN "11101000111" => data <= X"55000A58";
         WHEN "11101001000" => data <= X"6F6E6B6E";
         WHEN "11101001001" => data <= X"63206E77";
         WHEN "11101001010" => data <= X"2165646F";
         WHEN "11101001011" => data <= X"6F6E4B00";
         WHEN "11101001100" => data <= X"52206E77";
         WHEN "11101001101" => data <= X"32333253";
         WHEN "11101001110" => data <= X"6D6F6320";
         WHEN "11101001111" => data <= X"646E616D";
         WHEN "11101010000" => data <= X"000A3A73";
         WHEN "11101010001" => data <= X"53202A2A";
         WHEN "11101010010" => data <= X"74726174";
         WHEN "11101010011" => data <= X"65687420";
         WHEN "11101010100" => data <= X"6F727020";
         WHEN "11101010101" => data <= X"6D617267";
         WHEN "11101010110" => data <= X"616F6C20";
         WHEN "11101010111" => data <= X"20646564";
         WHEN "11101011000" => data <= X"74206E69";
         WHEN "11101011001" => data <= X"65677261";
         WHEN "11101011010" => data <= X"2A000A74";
         WHEN "11101011011" => data <= X"65532070";
         WHEN "11101011100" => data <= X"72702074";
         WHEN "11101011101" => data <= X"6172676F";
         WHEN "11101011110" => data <= X"6E696D6D";
         WHEN "11101011111" => data <= X"6F6D2067";
         WHEN "11101100000" => data <= X"28206564";
         WHEN "11101100001" => data <= X"61666564";
         WHEN "11101100010" => data <= X"29746C75";
         WHEN "11101100011" => data <= X"762A000A";
         WHEN "11101100100" => data <= X"74655320";
         WHEN "11101100101" => data <= X"72657620";
         WHEN "11101100110" => data <= X"63696669";
         WHEN "11101100111" => data <= X"6F697461";
         WHEN "11101101000" => data <= X"6F6D206E";
         WHEN "11101101001" => data <= X"000A6564";
         WHEN "11101101010" => data <= X"5320692A";
         WHEN "11101101011" => data <= X"20776F68";
         WHEN "11101101100" => data <= X"6F666E69";
         WHEN "11101101101" => data <= X"206E6F20";
         WHEN "11101101110" => data <= X"676F7270";
         WHEN "11101101111" => data <= X"206D6172";
         WHEN "11101110000" => data <= X"74206E69";
         WHEN "11101110001" => data <= X"65677261";
         WHEN "11101110010" => data <= X"2A000A74";
         WHEN "11101110011" => data <= X"6F542074";
         WHEN "11101110100" => data <= X"656C6767";
         WHEN "11101110101" => data <= X"72617420";
         WHEN "11101110110" => data <= X"20746567";
         WHEN "11101110111" => data <= X"77746562";
         WHEN "11101111000" => data <= X"206E6565";
         WHEN "11101111001" => data <= X"61524453";
         WHEN "11101111010" => data <= X"6428206D";
         WHEN "11101111011" => data <= X"75616665";
         WHEN "11101111100" => data <= X"2029746C";
         WHEN "11101111101" => data <= X"20646E61";
         WHEN "11101111110" => data <= X"73616C46";
         WHEN "11101111111" => data <= X"2A000A68";
         WHEN "11110000000" => data <= X"6550206D";
         WHEN "11110000001" => data <= X"726F6672";
         WHEN "11110000010" => data <= X"6973206D";
         WHEN "11110000011" => data <= X"656C706D";
         WHEN "11110000100" => data <= X"52445320";
         WHEN "11110000101" => data <= X"6D206D61";
         WHEN "11110000110" => data <= X"68636D65";
         WHEN "11110000111" => data <= X"0A6B6365";
         WHEN "11110001000" => data <= X"20732A00";
         WHEN "11110001001" => data <= X"63656843";
         WHEN "11110001010" => data <= X"5053206B";
         WHEN "11110001011" => data <= X"6C662D49";
         WHEN "11110001100" => data <= X"20687361";
         WHEN "11110001101" => data <= X"70696863";
         WHEN "11110001110" => data <= X"652A000A";
         WHEN "11110001111" => data <= X"61724520";
         WHEN "11110010000" => data <= X"53206573";
         WHEN "11110010001" => data <= X"662D4950";
         WHEN "11110010010" => data <= X"6873616C";
         WHEN "11110010011" => data <= X"69686320";
         WHEN "11110010100" => data <= X"2A000A70";
         WHEN "11110010101" => data <= X"75522072";
         WHEN "11110010110" => data <= X"7270206E";
         WHEN "11110010111" => data <= X"6172676F";
         WHEN "11110011000" => data <= X"6E69206D";
         WHEN "11110011001" => data <= X"49505320";
         WHEN "11110011010" => data <= X"616C662D";
         WHEN "11110011011" => data <= X"000A6873";
         WHEN "11110011100" => data <= X"5320662A";
         WHEN "11110011101" => data <= X"65726F74";
         WHEN "11110011110" => data <= X"6F727020";
         WHEN "11110011111" => data <= X"6D617267";
         WHEN "11110100000" => data <= X"616F6C20";
         WHEN "11110100001" => data <= X"20646564";
         WHEN "11110100010" => data <= X"53206E69";
         WHEN "11110100011" => data <= X"4D415244";
         WHEN "11110100100" => data <= X"206F7420";
         WHEN "11110100101" => data <= X"2D495053";
         WHEN "11110100110" => data <= X"73616C46";
         WHEN "11110100111" => data <= X"2A000A68";
         WHEN "11110101000" => data <= X"6F432063";
         WHEN "11110101001" => data <= X"7261706D";
         WHEN "11110101010" => data <= X"72702065";
         WHEN "11110101011" => data <= X"6172676F";
         WHEN "11110101100" => data <= X"6F6C206D";
         WHEN "11110101101" => data <= X"64656461";
         WHEN "11110101110" => data <= X"206E6920";
         WHEN "11110101111" => data <= X"41524453";
         WHEN "11110110000" => data <= X"6977204D";
         WHEN "11110110001" => data <= X"53206874";
         WHEN "11110110010" => data <= X"462D4950";
         WHEN "11110110011" => data <= X"6873616C";
         WHEN "11110110100" => data <= X"682A000A";
         WHEN "11110110101" => data <= X"69685420";
         WHEN "11110110110" => data <= X"65682073";
         WHEN "11110110111" => data <= X"6373706C";
         WHEN "11110111000" => data <= X"6E656572";
         WHEN "11110111001" => data <= X"00000A0A";
         WHEN "11110111010" => data <= X"EFBEADDE";
         WHEN "11110111011" => data <= X"01000000";
         WHEN "11110111100" => data <= X"02000000";
         WHEN "11110111101" => data <= X"03000000";
         WHEN "11110111110" => data <= X"04000000";
         WHEN "11110111111" => data <= X"05000000";
         WHEN "11111000000" => data <= X"06000000";
         WHEN "11111000001" => data <= X"07000000";
         WHEN "11111000010" => data <= X"2D1D00F0";
         WHEN "11111000011" => data <= X"441D00F0";
         WHEN "11111000100" => data <= X"6B1D00F0";
         WHEN "11111000101" => data <= X"8E1D00F0";
         WHEN "11111000110" => data <= X"A81D00F0";
         WHEN "11111000111" => data <= X"CB1D00F0";
         WHEN "11111001000" => data <= X"FF1D00F0";
         WHEN "11111001001" => data <= X"211E00F0";
         WHEN "11111001010" => data <= X"3A1E00F0";
         WHEN "11111001011" => data <= X"531E00F0";
         WHEN "11111001100" => data <= X"701E00F0";
         WHEN "11111001101" => data <= X"9F1E00F0";
         WHEN "11111001110" => data <= X"D21E00F0";
         WHEN "11111010000" => data <= X"10000000";
         WHEN "11111010010" => data <= X"00527A01";
         WHEN "11111010011" => data <= X"01097C04";
         WHEN "11111010100" => data <= X"00010D1B";
         WHEN "11111010101" => data <= X"14000000";
         WHEN "11111010110" => data <= X"18000000";
         WHEN "11111010111" => data <= X"64F8FFFF";
         WHEN "11111011000" => data <= X"14000000";
         WHEN "11111011001" => data <= X"09094100";
         WHEN "11111011010" => data <= X"0000000D";
         WHEN OTHERS => data <= X"00000000";
      END CASE;
   END PROCESS TheRom;

END platform_independent;
