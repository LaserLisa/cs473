../sandbox/bios_rom-behavior.vhdl